[32] filter_l [120][300][4] = {{{32'd2492, 32'd4439, 32'd6575, -32'd1302},
{-32'd9507, -32'd5766, -32'd8938, 32'd2714},
{32'd3401, 32'd9569, -32'd2886, 32'd9698},
{-32'd9913, 32'd8638, -32'd15976, 32'd3827},
{32'd8076, -32'd13545, -32'd8463, -32'd2571},
{-32'd314, -32'd1221, 32'd2466, 32'd15451},
{32'd7485, -32'd6844, -32'd8795, -32'd8492},
{32'd3171, -32'd10785, -32'd842, 32'd10965},
{32'd8588, 32'd8338, -32'd1251, 32'd4296},
{32'd5327, 32'd12892, 32'd2723, 32'd938},
{-32'd2901, -32'd3799, 32'd7386, 32'd1842},
{-32'd14012, -32'd109, 32'd4382, -32'd8304},
{32'd1700, 32'd4729, -32'd11259, 32'd3520},
{-32'd13295, -32'd10045, -32'd3068, -32'd1768},
{32'd484, -32'd7758, -32'd8764, -32'd2464},
{32'd1574, 32'd3251, -32'd10583, -32'd6721},
{-32'd147, -32'd374, 32'd7089, 32'd2154},
{32'd366, -32'd344, -32'd236, 32'd5896},
{-32'd2676, -32'd7507, -32'd3911, -32'd6968},
{32'd2037, -32'd4615, -32'd5722, -32'd4265},
{-32'd5011, 32'd5434, -32'd6266, 32'd5977},
{-32'd3081, -32'd3413, -32'd6431, -32'd4211},
{-32'd12694, -32'd796, -32'd3752, 32'd12845},
{32'd12399, -32'd9116, 32'd1663, -32'd5635},
{-32'd2455, 32'd10208, -32'd4850, 32'd1514},
{32'd7549, -32'd9267, 32'd2804, 32'd1013},
{32'd26, 32'd4372, -32'd7107, 32'd6545},
{-32'd3599, 32'd4821, -32'd9820, -32'd5444},
{-32'd1259, -32'd1317, -32'd8011, 32'd6361},
{32'd6771, 32'd1199, 32'd2579, -32'd3540},
{-32'd19547, 32'd8242, -32'd9770, 32'd7571},
{-32'd9017, -32'd12843, -32'd8251, 32'd2691},
{-32'd693, 32'd3104, 32'd14023, -32'd378},
{32'd2307, -32'd4258, -32'd2776, -32'd10533},
{32'd3657, 32'd7324, -32'd1241, 32'd1677},
{32'd19133, 32'd7936, 32'd3497, -32'd6248},
{-32'd2923, -32'd3644, 32'd4515, 32'd4408},
{-32'd8537, 32'd294, -32'd12511, -32'd6994},
{-32'd9053, -32'd5613, 32'd4058, 32'd2886},
{32'd12454, -32'd7465, 32'd13467, -32'd2859},
{32'd9276, 32'd12546, -32'd6625, -32'd12336},
{32'd12264, -32'd5103, -32'd8781, -32'd820},
{32'd1396, -32'd2011, -32'd9668, -32'd9605},
{-32'd1567, -32'd7849, -32'd1304, -32'd4592},
{32'd3045, -32'd4736, -32'd5803, -32'd1836},
{32'd6702, -32'd4753, 32'd4206, 32'd6820},
{-32'd10008, -32'd621, -32'd15059, -32'd6918},
{-32'd2394, -32'd8120, 32'd2575, 32'd10666},
{32'd7479, 32'd4110, -32'd15631, 32'd1731},
{-32'd12879, -32'd6525, -32'd6522, 32'd163},
{-32'd11604, 32'd774, 32'd3455, 32'd8286},
{-32'd1749, -32'd607, -32'd4513, -32'd15031},
{-32'd12166, -32'd9218, 32'd6009, 32'd4843},
{32'd1289, 32'd5973, 32'd7429, -32'd8255},
{32'd4667, 32'd949, 32'd6963, -32'd2821},
{-32'd5003, 32'd2191, 32'd397, 32'd4424},
{-32'd6168, 32'd548, 32'd2841, 32'd14735},
{-32'd2055, -32'd5046, 32'd9655, 32'd3541},
{32'd338, -32'd5429, -32'd929, -32'd4611},
{-32'd4445, -32'd9600, -32'd3996, 32'd13525},
{32'd10887, -32'd4257, -32'd8131, 32'd6748},
{-32'd2602, 32'd3429, -32'd6324, 32'd1042},
{32'd8277, -32'd4030, -32'd8047, -32'd3802},
{32'd2736, 32'd4373, -32'd8666, 32'd13330},
{-32'd1904, -32'd939, 32'd9851, 32'd187},
{32'd5081, 32'd46, 32'd5651, 32'd3304},
{-32'd5178, -32'd1598, 32'd3197, 32'd4836},
{-32'd11927, -32'd8671, -32'd36, 32'd6452},
{-32'd3507, -32'd5370, -32'd3663, -32'd5237},
{32'd1040, -32'd6239, 32'd914, 32'd8359},
{32'd3904, -32'd4202, 32'd3557, -32'd7172},
{32'd13192, 32'd2981, 32'd5414, -32'd7778},
{32'd412, -32'd3625, -32'd7280, -32'd12735},
{-32'd2841, 32'd13302, -32'd9964, 32'd17735},
{32'd3321, 32'd1032, 32'd8200, 32'd6072},
{32'd226, -32'd1592, 32'd11578, -32'd10483},
{-32'd10159, -32'd4126, 32'd1160, 32'd15755},
{32'd5058, 32'd2330, -32'd7592, 32'd7811},
{32'd12799, -32'd1002, -32'd4589, 32'd3534},
{32'd8843, 32'd3279, 32'd9667, 32'd838},
{-32'd4121, 32'd2932, 32'd1093, 32'd6350},
{32'd1292, -32'd1091, 32'd10884, -32'd1795},
{-32'd6759, 32'd3710, 32'd12419, 32'd1196},
{32'd6248, -32'd1836, 32'd6677, -32'd4124},
{32'd41, -32'd6907, 32'd4698, -32'd13379},
{-32'd4082, -32'd7337, 32'd3600, -32'd3910},
{32'd8145, 32'd2705, 32'd6122, -32'd8054},
{-32'd3678, -32'd3100, -32'd8286, -32'd6365},
{-32'd7049, -32'd8320, 32'd2050, 32'd7018},
{-32'd4591, -32'd4402, -32'd1361, 32'd7575},
{32'd791, 32'd3563, -32'd4658, -32'd4614},
{-32'd279, -32'd4895, -32'd11842, 32'd6316},
{32'd1522, -32'd1261, -32'd5585, -32'd1341},
{-32'd8265, -32'd5122, -32'd222, 32'd5205},
{32'd2887, -32'd9799, -32'd2711, -32'd5004},
{-32'd8299, -32'd1012, -32'd6012, 32'd1439},
{-32'd167, 32'd12685, 32'd15999, -32'd5730},
{32'd7449, 32'd8143, -32'd974, 32'd2594},
{32'd12449, -32'd11646, -32'd9065, 32'd1748},
{32'd2194, 32'd8772, 32'd11367, -32'd1362},
{-32'd5081, 32'd453, 32'd3331, 32'd11132},
{32'd75, -32'd2571, -32'd393, 32'd3086},
{32'd2329, 32'd5907, 32'd14271, -32'd7079},
{-32'd8776, 32'd8805, 32'd5993, 32'd11027},
{32'd7090, 32'd12228, 32'd721, 32'd4493},
{32'd2679, -32'd712, -32'd2564, 32'd9506},
{-32'd3766, 32'd2611, -32'd11488, -32'd2023},
{-32'd12752, 32'd7083, 32'd1145, -32'd1220},
{32'd5893, 32'd10397, 32'd10783, 32'd4732},
{-32'd3857, 32'd84, -32'd7450, 32'd7985},
{-32'd7742, 32'd6554, 32'd15662, -32'd3681},
{32'd12614, 32'd1330, 32'd13673, -32'd5171},
{-32'd1780, 32'd1938, 32'd11535, -32'd4528},
{32'd4469, 32'd2007, 32'd2535, -32'd3315},
{32'd8100, 32'd453, 32'd8424, -32'd2444},
{32'd7788, 32'd2180, -32'd11951, -32'd5593},
{32'd1193, 32'd4027, 32'd3883, -32'd5050},
{-32'd4805, 32'd7609, -32'd4175, 32'd7864},
{32'd949, 32'd9067, 32'd8305, -32'd8778},
{-32'd3138, 32'd6353, 32'd2118, 32'd1592},
{-32'd3492, 32'd7213, -32'd415, -32'd3752},
{32'd2808, -32'd2427, -32'd347, -32'd4959},
{-32'd13393, 32'd854, -32'd5357, 32'd5620},
{-32'd290, 32'd8766, -32'd9709, 32'd2508},
{-32'd10697, -32'd1410, 32'd8402, 32'd4833},
{-32'd5713, -32'd2474, 32'd4104, 32'd11007},
{32'd2532, 32'd4325, 32'd1796, -32'd3531},
{32'd3207, -32'd4868, -32'd4087, -32'd8643},
{32'd4569, -32'd10317, 32'd1539, 32'd5386},
{-32'd7190, 32'd3637, -32'd17855, -32'd2336},
{32'd578, -32'd1644, -32'd5881, -32'd9254},
{-32'd718, -32'd12358, -32'd9525, -32'd9796},
{-32'd17148, 32'd88, -32'd9098, -32'd4530},
{-32'd8412, -32'd6972, -32'd10699, 32'd3058},
{-32'd7165, -32'd231, -32'd7411, -32'd3500},
{32'd6287, -32'd4780, -32'd2245, -32'd574},
{32'd3712, -32'd1370, 32'd1231, 32'd6629},
{-32'd16228, -32'd1650, -32'd3280, 32'd6368},
{-32'd7557, 32'd463, 32'd8039, -32'd1737},
{32'd1510, -32'd2358, -32'd5512, 32'd2465},
{-32'd9590, 32'd8924, 32'd7627, 32'd2383},
{32'd3565, -32'd9836, 32'd1056, 32'd5455},
{-32'd9487, -32'd6264, 32'd6925, -32'd7289},
{-32'd13436, -32'd9050, -32'd22321, 32'd3977},
{32'd11, 32'd5160, 32'd12815, 32'd7651},
{-32'd5819, 32'd3891, 32'd5751, 32'd8087},
{-32'd4601, -32'd13166, 32'd2239, 32'd157},
{32'd8055, -32'd2538, 32'd1187, -32'd8036},
{32'd7857, 32'd3644, -32'd6446, 32'd4103},
{32'd1037, -32'd4074, -32'd5927, -32'd3392},
{-32'd1585, -32'd15639, 32'd2061, -32'd6901},
{32'd624, 32'd1659, -32'd527, -32'd512},
{-32'd1434, 32'd10332, 32'd5693, -32'd8696},
{-32'd3046, 32'd11269, 32'd4591, 32'd11225},
{32'd120, 32'd4684, -32'd11561, -32'd6039},
{32'd7575, -32'd2046, 32'd1722, -32'd12673},
{-32'd1843, 32'd7954, -32'd376, -32'd1086},
{-32'd3938, -32'd9334, -32'd513, 32'd5531},
{-32'd4088, -32'd3110, -32'd8419, -32'd8543},
{32'd12161, 32'd3356, -32'd12749, -32'd2594},
{32'd1337, 32'd4557, 32'd5893, -32'd2199},
{-32'd1963, -32'd697, 32'd2450, 32'd8003},
{-32'd8480, 32'd8119, -32'd2575, 32'd4386},
{-32'd1330, -32'd1917, 32'd14701, -32'd8807},
{32'd2824, 32'd5987, 32'd7291, 32'd1663},
{32'd917, -32'd1379, -32'd7834, 32'd7477},
{32'd5397, -32'd995, -32'd3429, 32'd5857},
{-32'd1810, -32'd12371, -32'd3372, -32'd3321},
{32'd15465, -32'd11743, -32'd31, -32'd6859},
{32'd11344, -32'd11572, 32'd3925, 32'd4625},
{32'd9414, 32'd6581, -32'd7695, 32'd2438},
{-32'd3408, -32'd4869, -32'd10195, 32'd2701},
{32'd6963, 32'd3781, 32'd5079, -32'd3460},
{-32'd8872, -32'd9399, -32'd5877, 32'd658},
{-32'd855, 32'd4622, 32'd2396, -32'd5808},
{32'd181, 32'd8688, -32'd5639, 32'd633},
{32'd232, 32'd951, -32'd3613, 32'd5221},
{-32'd4269, -32'd7528, -32'd1798, -32'd409},
{32'd7695, 32'd6702, 32'd6123, -32'd10119},
{-32'd623, -32'd10445, 32'd8146, 32'd5054},
{32'd5003, -32'd4264, 32'd14359, -32'd5814},
{-32'd7305, 32'd2186, 32'd2754, -32'd6893},
{-32'd13075, -32'd7814, 32'd519, 32'd5902},
{32'd1812, -32'd5094, -32'd4858, -32'd6057},
{-32'd11585, 32'd5101, 32'd5484, 32'd9251},
{-32'd3453, 32'd8257, 32'd3220, -32'd2121},
{32'd335, 32'd1683, -32'd12482, 32'd4531},
{-32'd10205, 32'd4516, 32'd15455, -32'd1460},
{32'd88, 32'd5671, -32'd1536, 32'd9661},
{-32'd1517, -32'd2078, -32'd6224, -32'd6812},
{32'd12648, -32'd4056, -32'd3468, -32'd7182},
{-32'd743, -32'd9760, 32'd1089, 32'd1797},
{-32'd9373, -32'd4624, 32'd5996, -32'd299},
{-32'd2836, 32'd3803, -32'd9599, 32'd19693},
{32'd975, -32'd5602, 32'd10238, 32'd295},
{-32'd4259, 32'd6277, -32'd4682, 32'd3586},
{-32'd7045, 32'd6089, 32'd4152, 32'd2589},
{-32'd1130, 32'd8239, -32'd4026, 32'd7546},
{-32'd700, 32'd510, -32'd5614, 32'd10440},
{-32'd6078, 32'd2794, 32'd2082, -32'd7097},
{-32'd3037, -32'd7579, -32'd221, -32'd804},
{32'd1797, -32'd434, 32'd3574, -32'd1780},
{-32'd1781, 32'd7233, 32'd5633, -32'd6807},
{-32'd3605, 32'd4160, 32'd6531, 32'd318},
{-32'd13788, -32'd6100, 32'd5401, 32'd13218},
{32'd7534, -32'd2203, -32'd6542, -32'd1491},
{-32'd770, 32'd24704, 32'd6439, 32'd7904},
{-32'd9365, -32'd1223, 32'd8566, 32'd4730},
{32'd1628, 32'd637, 32'd949, 32'd2929},
{-32'd5870, 32'd6960, 32'd10744, -32'd7395},
{-32'd772, -32'd10010, 32'd906, 32'd2287},
{-32'd7385, 32'd103, 32'd2368, 32'd9645},
{32'd2740, -32'd4191, 32'd3057, -32'd6667},
{32'd12449, -32'd7338, 32'd5418, 32'd1836},
{-32'd9955, -32'd5263, 32'd503, 32'd203},
{32'd2620, -32'd9086, -32'd4628, 32'd6435},
{32'd12406, 32'd4051, -32'd7536, 32'd5453},
{-32'd4679, -32'd8134, -32'd2095, 32'd1320},
{32'd4960, -32'd6843, 32'd13365, 32'd9845},
{32'd8161, -32'd1212, -32'd885, -32'd2110},
{-32'd5783, 32'd3755, 32'd7298, 32'd193},
{32'd753, 32'd7779, -32'd2093, -32'd5760},
{32'd8838, -32'd2763, 32'd7850, 32'd3403},
{32'd7137, 32'd5924, 32'd2127, -32'd8044},
{-32'd4893, -32'd1906, 32'd2300, 32'd17099},
{32'd10898, -32'd10994, 32'd5225, 32'd2778},
{-32'd13025, 32'd2968, 32'd666, 32'd2873},
{32'd3081, -32'd19387, -32'd1618, 32'd9680},
{-32'd11963, -32'd8532, 32'd6902, -32'd4211},
{32'd3835, 32'd7321, 32'd9760, -32'd2025},
{32'd3940, 32'd9004, 32'd2611, -32'd4557},
{32'd1644, 32'd10226, -32'd11833, -32'd11687},
{32'd6240, 32'd9364, 32'd5973, 32'd7013},
{-32'd8755, -32'd4197, 32'd954, 32'd2327},
{-32'd745, -32'd6206, -32'd542, -32'd7281},
{-32'd2479, -32'd10929, -32'd12955, -32'd12354},
{-32'd4051, 32'd14032, 32'd197, 32'd1238},
{-32'd1176, 32'd2195, -32'd9518, -32'd2203},
{32'd2770, 32'd5364, 32'd9501, -32'd4960},
{32'd1371, -32'd3025, 32'd3869, -32'd4682},
{32'd16177, 32'd6531, -32'd6152, 32'd1352},
{32'd7131, -32'd5934, 32'd7046, 32'd4123},
{-32'd4160, -32'd1715, -32'd2203, 32'd11889},
{-32'd1729, -32'd1601, -32'd514, 32'd18560},
{-32'd1356, 32'd14126, 32'd9587, 32'd2654},
{32'd2449, -32'd10145, 32'd3895, -32'd4264},
{32'd5428, -32'd6287, -32'd8958, -32'd4226},
{-32'd10597, 32'd8594, -32'd578, 32'd12295},
{32'd13836, -32'd2877, 32'd12066, 32'd3859},
{32'd6444, 32'd10003, 32'd8783, 32'd9105},
{32'd45, 32'd10104, -32'd11624, 32'd8742},
{-32'd2970, 32'd4079, -32'd5986, -32'd7109},
{-32'd1853, 32'd5390, 32'd675, -32'd2655},
{-32'd9456, 32'd360, 32'd11275, 32'd8933},
{32'd2135, 32'd4402, 32'd5577, -32'd10038},
{32'd14049, 32'd448, 32'd5342, -32'd5370},
{-32'd4171, 32'd4826, -32'd10909, -32'd201},
{-32'd9037, 32'd1446, -32'd2113, 32'd591},
{32'd7581, -32'd11623, -32'd1811, -32'd7242},
{32'd13613, -32'd400, 32'd11417, 32'd4734},
{-32'd1484, 32'd6094, -32'd15988, -32'd4215},
{32'd5765, -32'd6113, 32'd7052, -32'd13124},
{32'd4112, -32'd5687, 32'd8524, -32'd3930},
{32'd6818, -32'd421, 32'd5259, 32'd10427},
{-32'd12748, -32'd2195, 32'd2481, 32'd867},
{32'd3864, 32'd4823, 32'd20236, 32'd8366},
{32'd7068, -32'd8353, -32'd2560, -32'd3508},
{32'd2878, -32'd3423, -32'd4416, -32'd16846},
{32'd2255, -32'd16358, -32'd2770, -32'd10389},
{32'd1201, -32'd12910, 32'd4737, 32'd5069},
{32'd5329, -32'd11100, -32'd9498, 32'd15672},
{-32'd6075, 32'd261, -32'd5322, 32'd2149},
{32'd4575, -32'd3229, -32'd1954, -32'd10043},
{32'd2044, 32'd1621, 32'd4290, 32'd6902},
{-32'd10290, 32'd2610, 32'd6583, 32'd2076},
{-32'd818, -32'd6059, -32'd1813, 32'd2439},
{32'd5959, 32'd11840, 32'd5595, 32'd4366},
{32'd6588, -32'd2490, 32'd9075, -32'd2516},
{32'd146, -32'd7842, 32'd2446, -32'd1116},
{32'd1633, 32'd1160, -32'd6486, 32'd5257},
{-32'd1016, 32'd7248, -32'd2723, 32'd2043},
{-32'd1976, -32'd2840, -32'd2373, 32'd91},
{32'd4271, 32'd5780, -32'd14271, 32'd4718},
{32'd10512, -32'd2965, 32'd4072, 32'd11647},
{-32'd2501, 32'd10903, 32'd6566, -32'd2437},
{-32'd9387, -32'd6462, -32'd14783, 32'd2603},
{-32'd1491, 32'd353, -32'd8411, 32'd3620},
{32'd4896, -32'd923, -32'd7364, 32'd1775},
{32'd11379, -32'd13163, 32'd9166, 32'd1745},
{32'd8259, 32'd4120, -32'd247, -32'd8558},
{32'd11003, 32'd4086, -32'd549, -32'd7412},
{-32'd12609, 32'd9373, 32'd2530, 32'd10215},
{32'd1638, 32'd1646, -32'd4483, 32'd8338},
{-32'd1527, -32'd592, 32'd11909, 32'd4606},
{32'd4264, -32'd7513, -32'd6682, -32'd5388},
{32'd3272, -32'd12848, 32'd10660, -32'd6524},
{-32'd7077, 32'd5474, -32'd3466, -32'd6399},
{32'd12395, 32'd11086, 32'd4228, -32'd8225},
{-32'd2858, 32'd3511, -32'd4162, 32'd8105},
{32'd390, -32'd10642, 32'd1034, -32'd14110}
},
{{-32'd232, 32'd4849, 32'd5687, 32'd8795},
{-32'd7684, -32'd11861, -32'd9032, -32'd10620},
{32'd2663, -32'd3498, -32'd6092, 32'd8345},
{-32'd6120, 32'd9150, 32'd14020, 32'd3547},
{-32'd2004, -32'd11546, -32'd7064, -32'd9677},
{-32'd1006, 32'd6148, 32'd5776, -32'd4388},
{-32'd15895, -32'd10874, -32'd3466, 32'd2103},
{-32'd3216, -32'd6453, -32'd12940, -32'd6486},
{32'd7280, -32'd2144, 32'd5133, 32'd11248},
{32'd3612, 32'd15342, 32'd7954, 32'd13426},
{-32'd2028, 32'd7890, -32'd773, -32'd10057},
{-32'd310, 32'd6422, 32'd1583, -32'd4090},
{-32'd8244, 32'd13339, 32'd4357, -32'd2281},
{-32'd1930, -32'd11097, 32'd1134, 32'd5463},
{-32'd1417, -32'd4070, 32'd4122, -32'd5587},
{-32'd4019, -32'd6881, -32'd6396, -32'd2750},
{-32'd10192, 32'd13247, 32'd5521, 32'd5167},
{32'd6303, -32'd3576, -32'd8210, -32'd3550},
{32'd2919, -32'd3285, 32'd11798, 32'd3176},
{32'd4246, 32'd4504, -32'd2087, 32'd1849},
{32'd3568, -32'd2363, 32'd5369, -32'd20116},
{32'd6863, -32'd9800, 32'd9913, -32'd10484},
{-32'd8075, -32'd12728, -32'd3110, 32'd198},
{32'd415, 32'd470, -32'd6056, -32'd409},
{-32'd2767, 32'd8979, -32'd2933, 32'd5729},
{-32'd9683, 32'd6849, 32'd2312, -32'd4460},
{-32'd12527, -32'd12423, 32'd359, 32'd2327},
{32'd555, -32'd12479, 32'd4052, -32'd113},
{-32'd9766, -32'd1247, -32'd671, -32'd4889},
{32'd1907, -32'd6684, -32'd9707, -32'd3776},
{-32'd9005, 32'd17820, 32'd3359, 32'd5632},
{-32'd112, -32'd11845, -32'd8454, -32'd5566},
{-32'd9928, -32'd1487, 32'd6924, 32'd5458},
{-32'd190, -32'd8686, -32'd9985, -32'd9503},
{32'd3813, 32'd14503, -32'd990, 32'd11616},
{32'd15649, -32'd2576, -32'd4318, 32'd9914},
{32'd6452, -32'd10984, 32'd6282, 32'd9032},
{-32'd16086, 32'd18570, 32'd12023, 32'd1763},
{-32'd13411, 32'd8559, -32'd942, 32'd4234},
{-32'd4357, 32'd17653, -32'd4475, 32'd462},
{32'd756, -32'd3167, -32'd3, -32'd4309},
{32'd8521, -32'd6977, -32'd7918, 32'd1103},
{32'd909, 32'd6618, -32'd8819, -32'd6139},
{-32'd11410, -32'd78, -32'd5361, -32'd2954},
{32'd3280, 32'd3848, -32'd3008, -32'd4967},
{-32'd7999, -32'd10713, 32'd12563, 32'd4002},
{32'd1480, 32'd1475, -32'd1784, -32'd4914},
{-32'd7805, -32'd8386, 32'd5012, -32'd5769},
{32'd10880, 32'd2198, -32'd2849, 32'd3993},
{-32'd839, -32'd1070, -32'd12900, -32'd7074},
{-32'd6076, -32'd679, 32'd717, 32'd4314},
{32'd9570, -32'd4617, -32'd7025, 32'd639},
{32'd12677, -32'd6847, -32'd6880, -32'd17919},
{32'd10575, 32'd610, -32'd4444, 32'd1294},
{-32'd7125, 32'd64, -32'd5699, -32'd2009},
{-32'd1640, -32'd2593, 32'd12597, 32'd2104},
{-32'd8335, 32'd2596, 32'd1885, 32'd9522},
{-32'd8445, -32'd17832, 32'd3519, -32'd2927},
{32'd8684, -32'd4857, -32'd6702, -32'd1999},
{-32'd121, 32'd8380, -32'd2108, 32'd12776},
{32'd3941, -32'd18931, 32'd13967, 32'd2328},
{-32'd6641, -32'd728, 32'd4798, -32'd4249},
{32'd7711, 32'd382, -32'd2624, -32'd2537},
{32'd11943, -32'd3546, 32'd9033, 32'd138},
{-32'd5134, 32'd12146, 32'd4058, -32'd13482},
{-32'd6604, 32'd9479, 32'd2226, 32'd9250},
{-32'd6488, -32'd10153, 32'd11511, -32'd4534},
{32'd5608, -32'd3508, -32'd8378, -32'd10940},
{-32'd946, 32'd7197, -32'd3188, 32'd2141},
{32'd6329, 32'd3221, 32'd2525, -32'd844},
{-32'd14397, -32'd4513, 32'd9213, -32'd5452},
{-32'd20564, 32'd1877, -32'd12255, 32'd4967},
{32'd4572, -32'd7269, -32'd15437, 32'd11498},
{-32'd4682, -32'd676, -32'd5028, -32'd7472},
{-32'd9656, 32'd3624, 32'd13672, 32'd10534},
{-32'd4261, 32'd9047, -32'd1322, 32'd12753},
{-32'd4916, -32'd6055, -32'd8915, -32'd16273},
{-32'd10378, -32'd12443, -32'd380, -32'd1461},
{32'd2368, -32'd4997, 32'd4944, 32'd10009},
{32'd4301, -32'd3426, 32'd2491, 32'd6794},
{-32'd8060, -32'd10775, -32'd1843, -32'd1991},
{32'd1227, -32'd5081, -32'd5164, -32'd1606},
{32'd685, -32'd13966, 32'd10010, -32'd1533},
{32'd2003, 32'd4164, -32'd4602, -32'd4120},
{-32'd4360, 32'd4222, -32'd1953, -32'd12702},
{32'd5430, 32'd960, -32'd10531, -32'd4519},
{32'd8544, 32'd3593, -32'd340, 32'd12676},
{32'd3611, -32'd4325, 32'd5839, -32'd2973},
{-32'd6500, -32'd20873, 32'd7297, 32'd994},
{-32'd528, 32'd2991, 32'd5000, -32'd9565},
{-32'd3780, 32'd4700, -32'd7328, 32'd5258},
{-32'd6750, -32'd328, 32'd7051, -32'd12835},
{-32'd2188, 32'd7229, -32'd3145, 32'd315},
{32'd4772, -32'd5114, -32'd20524, -32'd2183},
{32'd5094, -32'd7440, -32'd7956, 32'd8991},
{-32'd5377, 32'd466, -32'd13606, -32'd16609},
{-32'd8938, 32'd6114, 32'd837, 32'd5658},
{32'd9364, 32'd3783, 32'd1595, 32'd4986},
{32'd3728, -32'd16163, -32'd780, -32'd7436},
{-32'd2033, 32'd6739, 32'd7923, 32'd7887},
{32'd4646, -32'd1717, -32'd4603, -32'd11529},
{32'd3466, 32'd3435, -32'd22655, 32'd1190},
{32'd3029, 32'd1928, 32'd2625, -32'd7558},
{-32'd94, 32'd21088, 32'd12440, 32'd7473},
{-32'd1193, 32'd10495, -32'd9600, 32'd1463},
{32'd7482, 32'd2246, -32'd1978, -32'd3975},
{32'd10715, -32'd6868, -32'd11771, 32'd631},
{-32'd10860, 32'd1003, -32'd14260, -32'd9511},
{-32'd5539, 32'd11347, -32'd2260, -32'd4455},
{32'd4732, 32'd2796, -32'd5161, 32'd4296},
{-32'd13036, -32'd13490, 32'd9693, -32'd1600},
{32'd9716, -32'd901, -32'd6349, 32'd3920},
{-32'd7979, 32'd12122, 32'd15603, 32'd4947},
{-32'd3640, -32'd16937, -32'd2532, -32'd9663},
{32'd3517, -32'd576, -32'd8779, 32'd2569},
{32'd5066, -32'd10583, -32'd4596, -32'd1714},
{32'd6693, 32'd10356, -32'd3638, -32'd2257},
{-32'd7429, 32'd669, -32'd15322, -32'd3050},
{-32'd7244, -32'd10071, -32'd7398, -32'd2552},
{32'd11470, 32'd7429, 32'd3337, 32'd8109},
{32'd2499, 32'd3143, -32'd15014, -32'd8652},
{32'd11786, -32'd2870, 32'd6590, 32'd7792},
{-32'd10300, -32'd11094, -32'd11207, -32'd9742},
{-32'd2554, 32'd4133, -32'd13597, -32'd40},
{32'd94, -32'd7101, 32'd6388, -32'd9722},
{-32'd643, 32'd17371, 32'd597, -32'd17},
{32'd4530, -32'd35, 32'd1306, -32'd5840},
{32'd1779, -32'd7481, 32'd655, -32'd1492},
{32'd5796, 32'd2342, -32'd11372, 32'd910},
{-32'd3036, -32'd9382, -32'd1988, -32'd2869},
{-32'd1503, 32'd1999, 32'd1940, 32'd8078},
{-32'd8878, 32'd5705, -32'd760, 32'd1610},
{32'd1694, -32'd916, 32'd2574, -32'd4029},
{-32'd5054, -32'd7290, -32'd10487, 32'd5436},
{-32'd2993, 32'd522, -32'd4054, 32'd3316},
{32'd3414, -32'd3041, -32'd3181, -32'd905},
{-32'd10590, -32'd17978, -32'd2740, 32'd2222},
{32'd7080, 32'd6745, 32'd2724, 32'd1466},
{32'd1266, -32'd1179, -32'd4479, 32'd3452},
{-32'd19880, -32'd16355, -32'd14359, -32'd3845},
{32'd3237, -32'd6229, -32'd4083, 32'd7625},
{-32'd3271, -32'd172, -32'd8410, -32'd2893},
{32'd5702, -32'd3415, -32'd8287, 32'd3160},
{-32'd10406, 32'd4406, -32'd2184, -32'd9204},
{32'd11395, 32'd4560, 32'd11159, 32'd8933},
{-32'd6590, -32'd11335, -32'd6114, 32'd4045},
{-32'd14726, 32'd2627, -32'd3318, -32'd11576},
{32'd1771, 32'd16159, 32'd16142, 32'd1541},
{-32'd1706, 32'd19399, 32'd10785, -32'd941},
{32'd7484, -32'd5241, -32'd1724, -32'd10017},
{-32'd6083, -32'd6531, -32'd4435, -32'd185},
{-32'd651, -32'd4319, 32'd3055, 32'd9054},
{-32'd85, 32'd1606, -32'd741, 32'd1615},
{32'd5585, 32'd607, -32'd1585, -32'd11866},
{-32'd7955, -32'd4930, -32'd7351, -32'd1261},
{-32'd2043, -32'd8346, 32'd7196, -32'd8731},
{32'd8600, 32'd4844, 32'd7317, 32'd15942},
{-32'd5073, 32'd7622, 32'd9590, -32'd1655},
{-32'd6941, -32'd13023, -32'd68, -32'd11328},
{32'd10448, 32'd10280, -32'd7227, 32'd1076},
{32'd12869, -32'd4906, -32'd9712, -32'd9554},
{32'd2935, -32'd8076, -32'd6624, 32'd9136},
{32'd757, -32'd2341, -32'd3752, -32'd4110},
{32'd4900, 32'd3905, -32'd6241, -32'd7873},
{32'd5043, 32'd17231, 32'd5772, 32'd9322},
{-32'd6828, 32'd9976, -32'd721, -32'd611},
{-32'd11779, 32'd314, -32'd1823, -32'd5718},
{-32'd3939, -32'd4747, 32'd5119, 32'd3423},
{-32'd4186, -32'd4179, -32'd1608, -32'd11191},
{32'd4150, 32'd4726, 32'd4908, -32'd6058},
{-32'd4816, -32'd7394, -32'd1259, -32'd9105},
{32'd17350, 32'd3255, 32'd6583, 32'd4104},
{32'd2568, 32'd16077, -32'd347, 32'd6344},
{-32'd1542, -32'd4, -32'd3121, -32'd8823},
{-32'd1515, 32'd1829, 32'd6631, -32'd1957},
{-32'd7521, 32'd11079, 32'd1168, -32'd2276},
{32'd4677, 32'd4031, 32'd8211, 32'd15101},
{-32'd6469, -32'd8313, 32'd2820, 32'd15818},
{32'd536, 32'd9907, 32'd1325, 32'd8066},
{-32'd6963, -32'd23715, 32'd6832, -32'd2926},
{-32'd2100, -32'd252, 32'd1452, 32'd221},
{-32'd8041, -32'd11764, -32'd8507, 32'd1362},
{32'd2315, -32'd5384, 32'd808, -32'd3144},
{-32'd6920, 32'd7665, -32'd185, -32'd7139},
{32'd11075, 32'd12938, -32'd9581, -32'd1009},
{-32'd206, 32'd1613, 32'd4540, 32'd930},
{32'd11626, 32'd5028, -32'd724, 32'd12128},
{-32'd14964, 32'd11193, -32'd16599, 32'd1874},
{-32'd12223, -32'd10211, -32'd8117, -32'd4591},
{32'd6726, -32'd13273, 32'd8476, 32'd2919},
{32'd10254, -32'd2351, -32'd15005, -32'd8289},
{-32'd10216, -32'd7241, -32'd9817, -32'd356},
{32'd3132, -32'd3390, -32'd1825, -32'd4667},
{32'd1744, -32'd12574, -32'd9925, 32'd6517},
{-32'd17838, -32'd6262, -32'd12396, 32'd4654},
{32'd2839, -32'd16361, 32'd250, -32'd9130},
{32'd10764, -32'd8835, 32'd2074, 32'd3085},
{-32'd2006, 32'd14150, 32'd9589, 32'd4466},
{-32'd6825, -32'd20615, 32'd4388, 32'd5169},
{-32'd5631, -32'd8809, -32'd11873, 32'd3673},
{32'd2634, -32'd11169, 32'd467, -32'd10127},
{-32'd1883, 32'd1291, -32'd19714, -32'd2380},
{-32'd3077, -32'd4683, -32'd5957, 32'd2769},
{-32'd4687, 32'd5022, 32'd12104, -32'd3135},
{-32'd4020, 32'd1674, 32'd3422, -32'd13279},
{-32'd3559, 32'd2048, -32'd5473, 32'd7806},
{32'd5518, 32'd9238, 32'd3114, -32'd2055},
{-32'd5468, -32'd312, 32'd753, -32'd15400},
{32'd371, -32'd12185, 32'd1362, 32'd15345},
{-32'd5144, -32'd4319, -32'd19694, -32'd7685},
{32'd854, -32'd7695, -32'd7088, -32'd1342},
{32'd3230, 32'd5224, 32'd606, 32'd1872},
{32'd32, 32'd2409, 32'd2740, -32'd11502},
{-32'd8795, 32'd1683, 32'd9838, -32'd1080},
{32'd3202, 32'd5144, 32'd2514, -32'd2222},
{-32'd363, -32'd3082, -32'd4374, 32'd3273},
{32'd10600, -32'd675, 32'd1005, 32'd4042},
{-32'd24561, -32'd3440, 32'd5449, 32'd3484},
{-32'd9586, 32'd12718, 32'd5827, 32'd7305},
{-32'd14956, 32'd1747, -32'd4798, -32'd2152},
{-32'd11227, -32'd2882, -32'd7410, -32'd2280},
{32'd4772, 32'd4144, 32'd7399, 32'd11861},
{-32'd2934, 32'd5749, -32'd8259, 32'd9943},
{-32'd1781, -32'd9386, -32'd7069, 32'd1098},
{32'd2231, -32'd9283, -32'd4440, -32'd6459},
{-32'd1867, -32'd3069, -32'd878, -32'd680},
{32'd917, 32'd2087, -32'd668, -32'd7148},
{32'd2178, -32'd24657, -32'd24177, 32'd1266},
{-32'd12865, -32'd3026, -32'd1399, 32'd9851},
{-32'd7968, 32'd1937, 32'd4402, 32'd7311},
{32'd8815, 32'd4343, -32'd10955, -32'd1733},
{-32'd2030, -32'd6900, 32'd576, 32'd3933},
{32'd10846, -32'd9917, 32'd9145, 32'd13366},
{32'd5000, -32'd2821, -32'd14178, -32'd4105},
{-32'd3138, -32'd5551, -32'd2505, -32'd1231},
{-32'd4153, -32'd14364, 32'd2681, -32'd4903},
{32'd73, 32'd5308, -32'd7094, -32'd3246},
{-32'd3409, 32'd1695, 32'd6378, 32'd5255},
{-32'd4900, -32'd7041, -32'd2468, 32'd7846},
{-32'd7865, -32'd9386, -32'd10218, -32'd4581},
{32'd8822, 32'd6886, 32'd4819, -32'd497},
{-32'd781, -32'd1149, 32'd7196, -32'd2371},
{-32'd4236, -32'd11495, -32'd5296, -32'd4233},
{32'd2224, 32'd2700, 32'd4731, 32'd7376},
{32'd1113, 32'd9902, 32'd1921, 32'd7423},
{32'd5565, -32'd7695, 32'd11011, 32'd319},
{-32'd12170, -32'd9869, -32'd10944, -32'd10249},
{32'd4895, -32'd2705, 32'd3076, -32'd13783},
{32'd607, 32'd8514, 32'd3532, -32'd180},
{-32'd5656, 32'd13461, 32'd14242, 32'd1618},
{32'd752, -32'd10663, -32'd5214, -32'd8246},
{32'd4175, -32'd2560, -32'd5438, -32'd9792},
{-32'd2259, -32'd493, 32'd8827, 32'd5320},
{-32'd5921, 32'd15528, 32'd3787, 32'd2439},
{-32'd7872, -32'd7121, -32'd16035, -32'd13907},
{32'd3452, -32'd797, 32'd8437, 32'd11643},
{-32'd2261, 32'd4139, 32'd5726, -32'd15724},
{-32'd5997, 32'd20953, 32'd9779, 32'd6528},
{32'd216, 32'd9302, -32'd4632, 32'd374},
{-32'd10628, 32'd43, -32'd3512, 32'd2886},
{32'd22792, 32'd4596, 32'd191, 32'd6167},
{32'd13681, -32'd13650, -32'd146, -32'd385},
{-32'd2467, -32'd4271, -32'd3296, 32'd651},
{32'd1685, -32'd9219, 32'd10270, 32'd12219},
{-32'd5454, 32'd9603, 32'd194, 32'd7588},
{32'd42, -32'd679, 32'd1572, 32'd7856},
{32'd10697, -32'd2701, 32'd7711, 32'd2951},
{32'd16708, -32'd5382, 32'd2567, 32'd8445},
{-32'd4518, 32'd4487, -32'd11021, -32'd6790},
{32'd2471, 32'd2237, 32'd16048, 32'd4748},
{-32'd2422, 32'd9729, 32'd5722, 32'd9348},
{-32'd1733, 32'd1950, 32'd4891, 32'd5054},
{-32'd9980, -32'd839, 32'd6183, -32'd14681},
{-32'd8752, 32'd5648, -32'd5612, 32'd965},
{-32'd7454, 32'd11916, -32'd3844, -32'd10911},
{-32'd2154, -32'd19041, 32'd8088, -32'd650},
{32'd5446, 32'd14370, 32'd7912, 32'd15310},
{-32'd487, -32'd1992, -32'd13581, -32'd8903},
{-32'd7855, -32'd11755, 32'd1264, -32'd3841},
{-32'd8408, -32'd4634, -32'd2228, 32'd2715},
{32'd17269, -32'd1259, -32'd2082, 32'd13396},
{-32'd2282, 32'd2377, 32'd9186, 32'd2784},
{-32'd4520, -32'd13623, -32'd6622, 32'd77},
{32'd5846, -32'd8287, 32'd4336, 32'd5146},
{-32'd13655, -32'd110, -32'd2047, 32'd11646},
{32'd109, -32'd6623, -32'd10207, -32'd9830},
{32'd11376, 32'd3009, 32'd13078, 32'd2647},
{32'd9920, -32'd3757, -32'd8713, -32'd6786},
{32'd744, 32'd8905, -32'd3342, 32'd1154},
{32'd2169, 32'd3240, -32'd6373, -32'd3926},
{-32'd2448, -32'd2835, 32'd10703, 32'd1239},
{32'd16164, 32'd15865, 32'd10765, 32'd5360},
{32'd3348, -32'd4841, 32'd10347, 32'd5601},
{32'd2211, -32'd3137, 32'd6368, -32'd8225},
{-32'd9671, 32'd4399, -32'd2080, -32'd2109},
{-32'd13958, -32'd10935, -32'd13880, -32'd6575},
{32'd6700, -32'd8076, -32'd5131, -32'd9578},
{32'd8017, 32'd9551, 32'd2674, 32'd5486},
{32'd6396, 32'd7614, 32'd3891, 32'd8683},
{32'd9251, 32'd1010, 32'd3722, 32'd6658}
},
{{-32'd4080, 32'd3846, 32'd10782, -32'd416},
{32'd1041, -32'd11186, 32'd1621, -32'd7696},
{32'd4053, -32'd10222, 32'd11076, 32'd1328},
{-32'd13005, 32'd6582, 32'd15810, 32'd13549},
{-32'd11419, 32'd2263, -32'd4724, 32'd8588},
{-32'd3343, -32'd541, 32'd1316, -32'd13495},
{-32'd1990, 32'd9737, -32'd7615, 32'd15901},
{32'd3697, -32'd7053, -32'd4791, -32'd6664},
{32'd6239, 32'd16060, 32'd2797, 32'd9279},
{-32'd9348, 32'd14977, 32'd10032, 32'd14610},
{32'd5323, -32'd14574, -32'd5741, -32'd1889},
{32'd6990, -32'd9051, 32'd973, 32'd8197},
{32'd925, -32'd2061, 32'd2765, -32'd5065},
{32'd4418, -32'd10196, -32'd1366, 32'd1277},
{32'd6873, -32'd3826, -32'd2167, 32'd2466},
{-32'd5213, 32'd919, -32'd10414, -32'd3031},
{-32'd4911, 32'd9299, 32'd12072, 32'd15343},
{32'd8646, 32'd5824, -32'd4185, 32'd1495},
{-32'd3792, 32'd1604, 32'd7807, 32'd1078},
{-32'd2119, 32'd8021, -32'd9995, -32'd2768},
{32'd10549, -32'd2817, 32'd1503, -32'd15599},
{-32'd6725, -32'd4154, 32'd5984, 32'd3011},
{32'd5431, 32'd5120, -32'd7165, 32'd8286},
{32'd13386, -32'd819, -32'd4693, -32'd8132},
{32'd2794, 32'd6213, 32'd6793, 32'd13042},
{32'd511, 32'd4251, 32'd9605, 32'd5050},
{-32'd1979, -32'd14943, 32'd3153, 32'd3517},
{-32'd3361, 32'd990, 32'd2354, -32'd5164},
{-32'd1349, 32'd5193, 32'd6401, -32'd740},
{-32'd665, -32'd8424, 32'd1754, -32'd8017},
{32'd580, 32'd14644, 32'd5326, 32'd10566},
{32'd13340, -32'd9156, -32'd6661, 32'd1040},
{-32'd15840, 32'd4238, 32'd12668, 32'd4357},
{32'd8027, -32'd13207, 32'd4459, -32'd1422},
{32'd2796, 32'd16591, 32'd6762, 32'd10106},
{32'd6142, -32'd4136, -32'd13710, 32'd4815},
{-32'd6371, 32'd4980, 32'd13454, 32'd414},
{-32'd15122, 32'd7574, 32'd4684, -32'd11101},
{-32'd8694, -32'd2891, -32'd7964, 32'd4164},
{-32'd7991, -32'd5545, -32'd9981, 32'd530},
{-32'd23632, 32'd3254, 32'd2546, -32'd7714},
{32'd12672, 32'd9548, -32'd10231, -32'd2692},
{-32'd1323, -32'd5479, 32'd3313, 32'd3791},
{32'd18724, -32'd6772, -32'd7096, -32'd3056},
{-32'd11064, -32'd10264, 32'd1802, 32'd15452},
{32'd3598, -32'd12343, -32'd4162, 32'd2946},
{32'd6988, -32'd3924, -32'd9816, -32'd4760},
{32'd10689, -32'd230, 32'd2814, -32'd10411},
{32'd1967, 32'd14414, -32'd9294, 32'd12329},
{32'd193, 32'd8269, -32'd1858, -32'd5051},
{-32'd2572, -32'd6537, -32'd10948, -32'd7692},
{-32'd2855, 32'd539, 32'd8590, 32'd7515},
{32'd14910, 32'd3412, -32'd11578, -32'd13004},
{32'd3718, -32'd6362, -32'd5753, 32'd4240},
{32'd1427, 32'd21245, -32'd2742, 32'd6018},
{-32'd11265, -32'd6018, 32'd8152, -32'd4865},
{-32'd96, 32'd8001, 32'd9258, -32'd155},
{-32'd11091, -32'd10724, -32'd16008, -32'd1150},
{32'd8665, 32'd2367, -32'd71, 32'd2139},
{32'd1431, 32'd703, -32'd2958, 32'd4710},
{32'd1457, -32'd5695, -32'd8827, 32'd11339},
{-32'd9518, 32'd3462, 32'd9637, -32'd3987},
{32'd3999, -32'd5814, -32'd10049, -32'd1698},
{-32'd709, 32'd3639, 32'd1444, 32'd1290},
{-32'd15835, -32'd1922, -32'd7444, 32'd6757},
{32'd15319, 32'd5466, 32'd4014, 32'd8898},
{-32'd5993, -32'd3406, 32'd7206, 32'd5918},
{32'd10230, 32'd6233, 32'd5908, -32'd7017},
{32'd4162, -32'd6164, 32'd1718, -32'd11183},
{32'd1619, 32'd863, -32'd2238, 32'd4987},
{32'd4291, -32'd4316, -32'd1134, -32'd2450},
{32'd7136, -32'd7522, 32'd6459, -32'd7077},
{32'd9333, -32'd8874, -32'd11721, -32'd566},
{32'd3360, 32'd4059, -32'd11548, 32'd3587},
{32'd7637, -32'd3049, 32'd10062, 32'd10449},
{32'd4698, 32'd5169, 32'd2594, -32'd2976},
{-32'd10759, -32'd1419, 32'd4650, -32'd6765},
{32'd4071, -32'd3044, 32'd5492, -32'd1430},
{32'd7067, 32'd12711, 32'd8412, -32'd5952},
{32'd5901, 32'd621, 32'd38, -32'd5723},
{-32'd4371, 32'd10704, -32'd5544, -32'd8183},
{-32'd7807, 32'd8277, 32'd1384, 32'd10993},
{-32'd4550, -32'd6847, -32'd17, 32'd3444},
{-32'd2336, 32'd7260, -32'd212, 32'd3324},
{32'd2562, 32'd6001, -32'd7683, -32'd7273},
{32'd8001, 32'd2000, 32'd5916, -32'd2967},
{-32'd10145, 32'd11116, 32'd411, 32'd485},
{-32'd8495, -32'd8682, -32'd13569, -32'd888},
{-32'd3200, -32'd3839, 32'd1989, -32'd9547},
{32'd3056, -32'd3419, 32'd1613, -32'd9749},
{-32'd6529, -32'd1405, -32'd1286, 32'd20926},
{32'd15544, -32'd7764, -32'd17003, -32'd8682},
{32'd2480, 32'd1185, 32'd3033, -32'd2599},
{32'd3578, 32'd9856, 32'd673, 32'd321},
{32'd13100, 32'd688, -32'd1072, -32'd1676},
{-32'd1789, -32'd704, -32'd1242, -32'd4260},
{-32'd10098, 32'd14591, 32'd11460, 32'd8918},
{32'd1461, 32'd1418, 32'd5077, -32'd212},
{32'd12507, -32'd2616, -32'd6229, -32'd3492},
{-32'd10872, 32'd15707, 32'd7753, 32'd10233},
{32'd17803, -32'd1983, 32'd8288, -32'd1989},
{-32'd3320, 32'd2364, -32'd3946, -32'd6720},
{32'd1627, 32'd6996, 32'd5272, 32'd9926},
{-32'd5958, -32'd1769, 32'd3232, 32'd853},
{-32'd9257, 32'd6921, 32'd1519, -32'd1208},
{32'd8978, -32'd869, -32'd5904, 32'd1648},
{32'd6059, -32'd15758, 32'd3427, -32'd4451},
{32'd20646, 32'd3573, 32'd3957, -32'd6596},
{-32'd1308, 32'd8256, -32'd3992, -32'd8765},
{32'd9006, -32'd4138, 32'd296, -32'd19160},
{32'd1901, -32'd5283, 32'd5183, -32'd6981},
{-32'd6249, 32'd1359, -32'd5959, 32'd10231},
{32'd4533, 32'd1784, 32'd1954, 32'd8952},
{-32'd6580, -32'd131, -32'd1510, 32'd23303},
{32'd3476, -32'd5340, -32'd83, -32'd7248},
{32'd9320, -32'd10009, -32'd8174, -32'd411},
{32'd10837, -32'd4912, -32'd841, 32'd9457},
{32'd4689, -32'd4924, 32'd963, -32'd1352},
{-32'd11568, -32'd15079, 32'd11272, 32'd7572},
{32'd10257, 32'd14564, 32'd351, 32'd1188},
{32'd14879, 32'd3052, -32'd5224, 32'd12632},
{-32'd2072, 32'd6412, 32'd13978, -32'd2685},
{-32'd6359, -32'd4025, 32'd1138, -32'd9357},
{-32'd825, -32'd10595, -32'd4479, 32'd4494},
{-32'd3004, 32'd3184, -32'd716, 32'd3582},
{32'd2203, 32'd10270, 32'd9683, -32'd11263},
{32'd650, -32'd3651, -32'd7080, -32'd5468},
{32'd7968, -32'd16025, 32'd604, -32'd9515},
{32'd663, -32'd8456, -32'd12953, -32'd11983},
{32'd5623, 32'd5645, -32'd764, 32'd5442},
{32'd9263, 32'd1435, -32'd19016, 32'd2744},
{-32'd5112, -32'd9214, -32'd2276, -32'd5673},
{-32'd6423, 32'd1563, -32'd1820, -32'd7026},
{-32'd383, -32'd10396, -32'd4390, -32'd2212},
{32'd8518, -32'd6568, 32'd5991, 32'd6041},
{32'd6245, -32'd1730, -32'd8908, -32'd354},
{32'd11797, -32'd3124, 32'd10010, -32'd6375},
{-32'd15170, -32'd938, 32'd2227, -32'd3170},
{32'd3368, 32'd3743, 32'd2094, -32'd2852},
{-32'd1090, 32'd547, -32'd5443, 32'd926},
{32'd849, -32'd6991, -32'd1231, -32'd5638},
{-32'd2863, -32'd10798, 32'd6053, -32'd3446},
{-32'd9747, -32'd671, 32'd2286, -32'd5136},
{-32'd804, 32'd6777, 32'd394, -32'd2473},
{32'd4435, -32'd2547, 32'd10457, 32'd9986},
{32'd3461, -32'd7634, 32'd5229, -32'd995},
{32'd17384, -32'd5660, -32'd820, -32'd7844},
{32'd5082, 32'd343, 32'd3536, 32'd4402},
{-32'd5913, 32'd541, 32'd8263, 32'd4396},
{-32'd8939, 32'd534, 32'd2416, 32'd1213},
{32'd689, -32'd5153, -32'd81, -32'd7875},
{-32'd10692, 32'd11845, 32'd3376, 32'd3234},
{-32'd5124, -32'd608, 32'd6994, -32'd1226},
{32'd4169, -32'd8240, -32'd226, 32'd8477},
{32'd10926, -32'd11144, -32'd2732, -32'd1320},
{-32'd1596, 32'd12395, 32'd1357, 32'd8807},
{32'd9096, 32'd3510, -32'd587, 32'd889},
{32'd21384, 32'd82, -32'd546, 32'd4271},
{-32'd4827, 32'd11199, 32'd4015, 32'd3493},
{-32'd4602, 32'd3554, 32'd337, 32'd3434},
{32'd8674, -32'd8361, -32'd16655, 32'd320},
{32'd1330, 32'd5432, 32'd15666, 32'd7225},
{32'd2293, -32'd14217, 32'd2724, -32'd3903},
{32'd4038, 32'd10070, 32'd12072, 32'd7114},
{32'd10968, 32'd104, 32'd172, -32'd5268},
{-32'd5500, 32'd848, -32'd9086, -32'd5592},
{32'd11013, -32'd4209, 32'd404, -32'd3107},
{-32'd1117, -32'd21251, -32'd4863, -32'd11805},
{-32'd8873, -32'd6817, 32'd1341, 32'd9708},
{32'd493, 32'd6015, -32'd12819, -32'd906},
{32'd3373, 32'd3084, 32'd2834, -32'd12834},
{32'd635, -32'd2554, -32'd695, -32'd7131},
{-32'd6314, 32'd11194, 32'd11591, 32'd10075},
{32'd3036, 32'd5512, -32'd9100, -32'd2439},
{32'd6984, -32'd4933, 32'd16129, 32'd2519},
{-32'd7253, -32'd4304, 32'd15351, -32'd4892},
{-32'd1962, 32'd3339, 32'd14161, 32'd8171},
{32'd1180, 32'd1387, -32'd3615, 32'd11290},
{32'd15877, 32'd5189, -32'd15090, 32'd1578},
{-32'd4347, -32'd18322, 32'd9477, -32'd408},
{32'd1548, 32'd5017, -32'd6253, 32'd4670},
{-32'd14140, 32'd5386, 32'd9760, -32'd4360},
{-32'd7426, -32'd7264, 32'd11211, -32'd6034},
{32'd5467, -32'd2743, 32'd4688, -32'd6832},
{32'd6872, -32'd8426, 32'd1199, -32'd1852},
{-32'd13896, 32'd13167, 32'd9005, 32'd711},
{32'd2749, -32'd1969, -32'd3239, 32'd1175},
{-32'd3081, 32'd9393, -32'd893, -32'd2325},
{32'd5240, 32'd843, -32'd8702, -32'd13929},
{-32'd11507, -32'd4559, -32'd1729, 32'd1659},
{-32'd7543, 32'd4875, -32'd10814, 32'd3669},
{32'd6732, -32'd8516, -32'd4710, -32'd7867},
{32'd7532, -32'd5369, -32'd2240, -32'd12086},
{32'd7768, -32'd5329, 32'd1713, -32'd1820},
{-32'd338, -32'd7811, 32'd3192, -32'd3731},
{-32'd4597, -32'd2183, 32'd1649, 32'd3299},
{-32'd4435, 32'd1407, 32'd9489, 32'd4936},
{-32'd6130, 32'd1419, 32'd6327, 32'd3113},
{-32'd12558, 32'd2110, -32'd2009, 32'd3345},
{-32'd1994, 32'd10016, -32'd2133, 32'd6888},
{32'd509, -32'd10070, -32'd9048, -32'd8986},
{32'd6626, -32'd7032, 32'd9252, -32'd9313},
{-32'd13784, -32'd716, -32'd6488, 32'd14095},
{-32'd7394, -32'd3978, -32'd5506, 32'd2157},
{32'd58, -32'd4560, -32'd2393, 32'd1343},
{-32'd4454, -32'd9707, 32'd5467, -32'd3063},
{-32'd6810, -32'd610, 32'd12577, 32'd4426},
{32'd10997, -32'd7827, -32'd3180, -32'd6403},
{32'd3095, 32'd9895, 32'd6172, -32'd7421},
{-32'd7632, 32'd802, 32'd14127, 32'd10608},
{-32'd2643, -32'd6135, 32'd3487, -32'd16601},
{32'd1514, -32'd1410, -32'd9840, 32'd1622},
{-32'd13623, -32'd545, -32'd512, -32'd1861},
{32'd7371, 32'd1363, 32'd2645, 32'd6925},
{32'd9349, 32'd606, 32'd2979, 32'd5011},
{32'd4631, -32'd2542, 32'd5079, -32'd9227},
{32'd5704, -32'd11809, -32'd1740, 32'd6438},
{32'd4735, -32'd5889, 32'd9538, -32'd11609},
{-32'd10128, 32'd7211, 32'd20586, 32'd3396},
{32'd9466, -32'd6054, 32'd3207, 32'd10865},
{32'd417, -32'd18236, -32'd1398, 32'd59},
{32'd12010, 32'd2886, -32'd732, 32'd11771},
{32'd8513, 32'd7409, -32'd10132, -32'd3351},
{32'd5021, 32'd4920, -32'd7874, -32'd3674},
{32'd6526, -32'd14574, -32'd5059, -32'd2269},
{32'd2499, -32'd4194, -32'd9165, 32'd10875},
{32'd11801, -32'd9546, -32'd2762, -32'd5701},
{-32'd2017, 32'd893, -32'd11548, -32'd4691},
{-32'd3239, -32'd6932, 32'd2763, -32'd5640},
{-32'd12418, -32'd7518, 32'd21806, 32'd4084},
{-32'd1908, -32'd9280, -32'd45, -32'd7066},
{-32'd1954, -32'd11550, -32'd9306, 32'd628},
{-32'd9035, 32'd11245, 32'd12790, 32'd1914},
{32'd2337, -32'd1636, 32'd1826, -32'd5071},
{-32'd9415, -32'd13206, -32'd4175, -32'd448},
{32'd10016, -32'd11106, -32'd2928, -32'd4553},
{-32'd9088, -32'd5756, -32'd7749, 32'd257},
{-32'd12468, 32'd1041, 32'd1216, -32'd847},
{-32'd6298, -32'd25, 32'd12104, 32'd536},
{-32'd265, 32'd2266, 32'd3005, 32'd8733},
{-32'd8843, -32'd3150, -32'd1144, -32'd4671},
{32'd292, -32'd895, 32'd5000, 32'd1265},
{-32'd2377, -32'd11213, -32'd7624, -32'd1839},
{-32'd5991, 32'd9210, -32'd1392, 32'd4162},
{-32'd7385, 32'd6033, 32'd13812, 32'd6592},
{-32'd3770, 32'd3543, 32'd12418, 32'd13965},
{-32'd6994, 32'd4556, 32'd1051, 32'd5507},
{32'd8111, 32'd164, -32'd3968, 32'd678},
{-32'd123, -32'd1793, 32'd5445, 32'd11166},
{-32'd1836, -32'd11556, 32'd6712, 32'd1660},
{32'd1223, -32'd1176, 32'd10449, -32'd13016},
{32'd6882, 32'd2241, -32'd3647, -32'd584},
{-32'd5835, 32'd5452, 32'd8697, 32'd12163},
{-32'd6114, -32'd1679, -32'd5936, -32'd363},
{-32'd3175, -32'd7310, -32'd7064, -32'd3217},
{-32'd647, -32'd486, -32'd1036, 32'd7685},
{-32'd7387, 32'd9499, -32'd7035, -32'd5601},
{-32'd5476, 32'd525, -32'd3816, 32'd486},
{-32'd7476, 32'd6651, -32'd11525, 32'd5886},
{32'd461, -32'd6984, 32'd6630, -32'd4495},
{32'd49, 32'd7895, -32'd1964, 32'd3175},
{32'd7726, -32'd3778, -32'd12260, -32'd2601},
{32'd1089, 32'd3951, -32'd1683, -32'd1427},
{32'd1162, -32'd9850, -32'd859, 32'd1623},
{32'd6198, 32'd9587, 32'd6378, -32'd6301},
{-32'd16554, 32'd11651, 32'd4075, 32'd5885},
{-32'd1024, 32'd10071, -32'd17351, -32'd3595},
{-32'd8907, 32'd7856, 32'd11575, 32'd10399},
{32'd17367, 32'd5659, -32'd15406, 32'd10500},
{-32'd2197, -32'd469, 32'd1475, -32'd2420},
{32'd15541, 32'd2323, 32'd9516, -32'd6054},
{32'd7200, 32'd3971, 32'd733, -32'd5252},
{-32'd6791, -32'd1771, -32'd716, -32'd18},
{32'd12502, -32'd8923, 32'd7497, -32'd13586},
{-32'd1931, 32'd3669, 32'd5441, -32'd6577},
{32'd8277, -32'd17565, -32'd820, -32'd7206},
{-32'd7061, 32'd19412, 32'd12402, 32'd13907},
{32'd10918, 32'd5002, -32'd12338, -32'd10407},
{32'd1895, -32'd8660, 32'd2056, -32'd2123},
{-32'd383, -32'd1618, 32'd201, -32'd2433},
{-32'd10693, 32'd3363, 32'd8462, 32'd9692},
{32'd2102, -32'd11505, -32'd12686, -32'd5714},
{32'd4167, 32'd9949, 32'd4880, 32'd7754},
{-32'd1696, -32'd7598, 32'd7833, -32'd7447},
{32'd5999, -32'd1574, 32'd3646, -32'd5686},
{-32'd12011, 32'd409, -32'd11843, 32'd3710},
{32'd556, 32'd7659, -32'd11404, -32'd4284},
{-32'd1986, 32'd5815, 32'd3072, -32'd11796},
{32'd4048, -32'd10249, -32'd11436, 32'd4264},
{32'd2238, 32'd2237, -32'd4506, 32'd3747},
{32'd12077, 32'd7870, -32'd8331, -32'd5772},
{32'd9534, 32'd3486, 32'd5170, 32'd8079},
{-32'd14988, 32'd15402, 32'd8573, 32'd1021},
{32'd632, 32'd2215, 32'd3505, -32'd3704},
{32'd1436, 32'd7377, -32'd1807, -32'd7138},
{32'd11138, -32'd3186, 32'd1389, -32'd8974},
{32'd2898, -32'd2995, -32'd5477, 32'd13989},
{-32'd7291, 32'd2729, 32'd2365, 32'd14915},
{32'd4897, 32'd12639, 32'd2850, -32'd2227},
{32'd10948, 32'd6555, -32'd5232, 32'd6945}
},
{{32'd8665, 32'd7787, -32'd2143, -32'd773},
{-32'd12248, 32'd1000, -32'd7542, 32'd598},
{-32'd4059, 32'd6364, 32'd7740, 32'd8333},
{-32'd5229, 32'd1729, 32'd13176, 32'd1624},
{32'd1678, 32'd4802, 32'd13011, 32'd22034},
{32'd2368, 32'd3531, -32'd1650, 32'd7304},
{32'd7970, -32'd3124, 32'd7626, -32'd2654},
{-32'd1414, -32'd252, -32'd3394, -32'd3090},
{32'd8313, 32'd3749, -32'd2885, 32'd4855},
{32'd321, 32'd5873, -32'd2041, -32'd4538},
{-32'd3360, -32'd4658, 32'd3939, 32'd10924},
{-32'd2501, -32'd3109, 32'd8996, -32'd2687},
{-32'd9522, -32'd15372, 32'd599, 32'd5711},
{32'd3444, 32'd826, 32'd388, -32'd9409},
{-32'd4913, 32'd2832, 32'd704, 32'd1561},
{32'd6046, -32'd465, 32'd8390, 32'd4749},
{32'd13164, 32'd1381, 32'd7053, 32'd6305},
{-32'd6361, -32'd517, -32'd3564, 32'd1847},
{32'd348, 32'd13185, -32'd7025, -32'd4674},
{32'd24442, 32'd6045, -32'd6758, 32'd7722},
{32'd3038, -32'd4040, -32'd9159, 32'd1456},
{32'd5116, -32'd12643, -32'd7484, -32'd6380},
{32'd1483, 32'd3134, -32'd8581, 32'd5175},
{-32'd7905, 32'd7512, 32'd11095, -32'd3140},
{-32'd1202, 32'd9055, -32'd1930, -32'd3844},
{-32'd4456, -32'd10020, 32'd19838, 32'd11146},
{-32'd1151, -32'd10459, -32'd10462, 32'd3445},
{-32'd5298, 32'd1846, -32'd2584, -32'd2262},
{32'd12119, 32'd7870, -32'd1280, -32'd8083},
{32'd10814, 32'd4547, -32'd2110, 32'd7899},
{32'd3120, 32'd11127, 32'd18018, 32'd7491},
{-32'd5170, -32'd9275, 32'd1820, -32'd1780},
{32'd3754, 32'd4745, 32'd9143, -32'd2694},
{32'd4522, -32'd6955, 32'd12407, 32'd98},
{-32'd2279, -32'd253, 32'd1268, -32'd1328},
{-32'd3019, 32'd2301, 32'd3687, -32'd5156},
{-32'd18775, 32'd11837, -32'd5662, -32'd7236},
{32'd5491, 32'd7481, -32'd99, -32'd2488},
{32'd3444, -32'd2062, -32'd2741, -32'd6478},
{32'd4447, -32'd11455, -32'd10057, 32'd11225},
{-32'd4718, -32'd2508, 32'd2574, -32'd3858},
{-32'd3750, -32'd6535, 32'd1685, 32'd2933},
{-32'd2066, 32'd9219, 32'd3435, 32'd8851},
{-32'd5439, -32'd3679, -32'd1188, 32'd6933},
{-32'd1704, 32'd2719, -32'd6947, -32'd14358},
{32'd3858, 32'd2229, -32'd6530, 32'd5130},
{-32'd2491, -32'd7326, -32'd14688, -32'd1692},
{-32'd6955, -32'd1911, 32'd8008, 32'd3473},
{-32'd8770, 32'd5566, -32'd9750, -32'd2943},
{-32'd8607, -32'd10449, -32'd5027, -32'd5846},
{32'd7385, -32'd10274, -32'd726, 32'd5664},
{32'd2791, -32'd578, -32'd3394, -32'd8933},
{-32'd7206, 32'd9981, 32'd5468, -32'd19523},
{-32'd4303, 32'd9715, 32'd13159, -32'd2270},
{-32'd3940, 32'd9019, 32'd3693, 32'd12188},
{32'd4294, -32'd12581, -32'd13129, -32'd109},
{32'd3339, -32'd10709, -32'd1916, 32'd1639},
{-32'd304, 32'd1941, 32'd924, -32'd651},
{-32'd1653, 32'd9900, -32'd8889, -32'd7592},
{32'd6371, -32'd7702, 32'd844, -32'd1755},
{-32'd634, -32'd11776, 32'd4262, 32'd18094},
{32'd896, 32'd3562, 32'd5039, 32'd720},
{-32'd8940, -32'd12624, 32'd3516, -32'd2867},
{-32'd6152, -32'd5659, -32'd1258, -32'd2621},
{-32'd1743, 32'd9621, -32'd13221, -32'd13303},
{32'd6251, -32'd2497, -32'd3974, -32'd8102},
{-32'd2526, 32'd4076, -32'd1492, 32'd9843},
{32'd2039, 32'd4577, 32'd3240, 32'd5560},
{-32'd3831, -32'd4265, -32'd4543, -32'd3857},
{32'd698, -32'd7195, 32'd2792, -32'd21269},
{32'd1645, 32'd5548, -32'd14206, 32'd7421},
{-32'd11894, -32'd3677, -32'd8189, 32'd408},
{-32'd15147, -32'd9283, -32'd3409, 32'd4284},
{32'd13180, -32'd7382, -32'd7371, -32'd9257},
{32'd12350, -32'd3249, 32'd6734, 32'd3753},
{-32'd4497, 32'd11324, 32'd8096, 32'd5922},
{-32'd1885, 32'd7265, -32'd4728, -32'd5144},
{32'd7503, 32'd2452, 32'd5590, -32'd4689},
{-32'd3837, 32'd4441, -32'd3129, -32'd2361},
{-32'd13830, -32'd2510, 32'd10200, 32'd4359},
{-32'd3139, 32'd15083, 32'd10826, -32'd3609},
{-32'd2948, -32'd7871, -32'd9536, -32'd14703},
{32'd5195, 32'd205, 32'd3150, 32'd423},
{32'd5425, -32'd997, 32'd2332, 32'd7767},
{32'd1942, -32'd12153, 32'd5552, 32'd2671},
{-32'd13936, -32'd728, -32'd2057, -32'd3047},
{-32'd4132, -32'd8142, -32'd200, -32'd1088},
{-32'd2722, 32'd2557, 32'd8344, 32'd335},
{32'd9067, 32'd6275, -32'd12581, -32'd12461},
{-32'd5266, -32'd2201, -32'd13622, -32'd7935},
{32'd2964, 32'd2939, -32'd3714, -32'd2393},
{32'd1991, -32'd17389, -32'd16763, -32'd3741},
{-32'd9200, 32'd17100, 32'd1754, -32'd2402},
{-32'd2538, 32'd10557, 32'd8488, 32'd10657},
{-32'd1114, 32'd208, 32'd3326, -32'd10795},
{-32'd10500, 32'd4386, -32'd4364, 32'd8914},
{32'd278, 32'd13697, 32'd15943, -32'd4607},
{-32'd6186, 32'd6733, 32'd19228, -32'd3305},
{-32'd1684, -32'd880, 32'd3087, -32'd1879},
{-32'd4114, 32'd7557, 32'd6679, -32'd1602},
{-32'd11, -32'd3304, 32'd2401, -32'd5359},
{32'd4156, 32'd15562, 32'd1006, -32'd11999},
{32'd3710, 32'd878, 32'd2011, 32'd4963},
{-32'd2320, -32'd1239, -32'd3421, 32'd1607},
{32'd1997, -32'd566, 32'd7469, 32'd2824},
{32'd2407, -32'd1563, -32'd3364, 32'd3511},
{-32'd8640, -32'd2450, 32'd9852, -32'd379},
{32'd5166, 32'd1488, 32'd11993, 32'd2742},
{-32'd4254, 32'd10273, -32'd6901, -32'd3274},
{-32'd1051, -32'd257, -32'd2585, 32'd1577},
{-32'd2163, -32'd2605, -32'd7915, 32'd1905},
{32'd4626, 32'd7231, -32'd10575, -32'd10276},
{32'd3456, 32'd1921, -32'd10925, -32'd11988},
{32'd5259, -32'd6046, 32'd3891, -32'd5603},
{-32'd2125, 32'd5567, 32'd1183, -32'd2599},
{32'd2580, 32'd452, -32'd14835, 32'd1944},
{32'd7864, 32'd840, 32'd4741, 32'd1236},
{32'd2876, 32'd9038, -32'd1240, 32'd2517},
{-32'd3033, -32'd8656, -32'd1290, -32'd4813},
{-32'd12159, -32'd6144, -32'd1174, -32'd300},
{-32'd6086, -32'd4799, -32'd7312, 32'd10458},
{-32'd7861, 32'd13337, 32'd13591, -32'd1634},
{-32'd3805, -32'd3737, 32'd1826, -32'd1348},
{32'd2397, -32'd4069, -32'd3302, -32'd1154},
{-32'd4324, -32'd12446, -32'd4287, 32'd17395},
{-32'd6017, 32'd5282, -32'd6991, 32'd2248},
{-32'd6426, -32'd2519, 32'd5184, 32'd2785},
{-32'd1975, -32'd466, -32'd5248, 32'd1900},
{-32'd7831, -32'd3892, -32'd860, 32'd18435},
{32'd3935, -32'd5395, 32'd16763, -32'd11042},
{32'd8176, -32'd10600, 32'd8934, 32'd12260},
{32'd11341, 32'd5899, 32'd515, -32'd4686},
{32'd2592, -32'd3842, 32'd1844, 32'd2448},
{-32'd933, -32'd1389, -32'd10345, -32'd807},
{32'd56, -32'd4669, 32'd1485, -32'd15659},
{-32'd2298, -32'd4748, -32'd5860, -32'd4625},
{32'd1048, -32'd4673, 32'd2482, 32'd2270},
{-32'd10276, 32'd11423, -32'd3407, -32'd4838},
{32'd3160, 32'd13376, 32'd4194, 32'd7732},
{-32'd3095, -32'd2543, -32'd11060, -32'd2020},
{-32'd5678, -32'd12171, 32'd6897, 32'd3509},
{32'd7212, -32'd11500, 32'd8966, 32'd1369},
{-32'd1612, -32'd1209, -32'd12053, 32'd342},
{-32'd2556, 32'd10919, 32'd8336, 32'd10861},
{-32'd955, 32'd1159, 32'd3086, 32'd2353},
{-32'd93, 32'd4647, 32'd440, 32'd5056},
{32'd7414, -32'd3398, -32'd1420, 32'd12339},
{-32'd417, -32'd6728, 32'd1698, 32'd5371},
{32'd1518, 32'd6424, 32'd8344, -32'd961},
{-32'd23411, -32'd9706, -32'd1339, 32'd4681},
{-32'd10824, 32'd9022, 32'd12539, 32'd7448},
{32'd7270, 32'd8042, -32'd5767, -32'd1580},
{32'd2344, -32'd7042, 32'd10777, 32'd4594},
{32'd1554, 32'd5496, 32'd3477, 32'd8992},
{-32'd4748, -32'd4513, -32'd9644, -32'd5609},
{-32'd5935, -32'd2351, 32'd6185, 32'd5394},
{32'd3258, -32'd6413, 32'd129, -32'd9456},
{32'd286, 32'd11443, -32'd2901, -32'd6260},
{32'd5028, 32'd5288, 32'd3583, -32'd6247},
{32'd2401, -32'd4031, -32'd3729, -32'd5479},
{-32'd2249, -32'd4361, -32'd6774, -32'd10286},
{-32'd5927, 32'd5654, 32'd9291, 32'd9515},
{32'd4542, -32'd3092, 32'd3129, -32'd11196},
{-32'd1677, 32'd3928, 32'd4773, -32'd11061},
{32'd13772, -32'd2274, -32'd11692, -32'd839},
{-32'd7770, -32'd6785, -32'd15224, -32'd6051},
{32'd8136, 32'd5446, 32'd6518, 32'd1259},
{32'd5979, -32'd11158, -32'd7210, -32'd173},
{-32'd4125, -32'd4658, 32'd7, 32'd5926},
{32'd6431, -32'd8633, 32'd10548, 32'd4510},
{-32'd6085, 32'd7241, -32'd6138, 32'd4317},
{-32'd1543, -32'd7537, 32'd7634, 32'd2503},
{32'd4252, -32'd3602, -32'd2251, 32'd973},
{-32'd11016, -32'd959, 32'd9096, -32'd6162},
{-32'd7696, -32'd2215, 32'd5262, -32'd7222},
{32'd9068, -32'd5, 32'd5085, -32'd3119},
{32'd3894, 32'd1513, 32'd12132, 32'd10310},
{32'd8342, 32'd12189, -32'd12419, -32'd3809},
{32'd5607, -32'd10516, 32'd1913, 32'd13650},
{-32'd4862, 32'd4219, 32'd1895, 32'd5451},
{32'd8721, -32'd4693, -32'd740, -32'd9501},
{-32'd6398, 32'd11990, 32'd3517, -32'd2639},
{-32'd4525, 32'd262, -32'd6685, -32'd6749},
{-32'd2681, 32'd6477, -32'd645, -32'd990},
{-32'd4167, -32'd3913, -32'd1386, 32'd6827},
{32'd12924, -32'd4427, -32'd172, 32'd1126},
{32'd745, 32'd1284, -32'd9061, -32'd4333},
{32'd2762, 32'd3833, 32'd419, -32'd10529},
{32'd10020, 32'd1783, -32'd13481, -32'd758},
{-32'd3772, -32'd1372, -32'd6353, -32'd9047},
{-32'd1191, -32'd1399, 32'd4424, 32'd718},
{-32'd5148, -32'd1005, -32'd7196, 32'd5152},
{-32'd9905, -32'd1529, -32'd13091, 32'd3409},
{-32'd12747, -32'd1688, -32'd7533, -32'd6033},
{32'd424, 32'd6021, -32'd2384, -32'd7838},
{-32'd1579, 32'd6848, 32'd4149, 32'd7820},
{-32'd10608, 32'd5019, 32'd1341, 32'd3610},
{32'd12483, -32'd2672, 32'd2438, -32'd3448},
{-32'd15060, -32'd910, -32'd4266, 32'd6074},
{32'd1249, 32'd16650, 32'd7027, 32'd8603},
{32'd535, -32'd1657, -32'd14067, 32'd3422},
{-32'd10521, -32'd855, 32'd14711, 32'd13614},
{32'd4370, -32'd5736, -32'd462, 32'd7519},
{-32'd7469, -32'd1507, -32'd6756, 32'd1801},
{32'd3186, -32'd3554, -32'd15628, -32'd6237},
{-32'd3908, -32'd9205, -32'd546, 32'd846},
{32'd9217, 32'd4329, 32'd9195, -32'd6658},
{32'd4132, -32'd5625, -32'd18898, -32'd12392},
{-32'd5754, 32'd2196, 32'd5440, 32'd9017},
{32'd611, 32'd14515, 32'd7529, 32'd2977},
{-32'd11912, 32'd194, 32'd927, 32'd11192},
{32'd1064, 32'd536, -32'd14132, -32'd2997},
{32'd1457, -32'd8178, -32'd4372, 32'd2643},
{-32'd5050, 32'd5829, -32'd72, -32'd5845},
{-32'd15039, 32'd3832, 32'd1297, 32'd14669},
{32'd2691, -32'd33, 32'd6975, -32'd706},
{32'd10166, 32'd2508, 32'd2511, -32'd2962},
{-32'd8525, -32'd936, -32'd2316, -32'd911},
{32'd13996, 32'd9268, 32'd8291, -32'd926},
{-32'd428, -32'd5538, 32'd2448, 32'd193},
{32'd15933, 32'd4873, 32'd6721, 32'd12923},
{32'd3044, -32'd9364, -32'd5391, 32'd2102},
{-32'd4316, 32'd15419, -32'd1398, 32'd4675},
{-32'd3501, -32'd4971, 32'd152, -32'd8037},
{32'd3722, -32'd2954, 32'd2430, 32'd657},
{-32'd2771, -32'd3689, -32'd542, -32'd5118},
{32'd14269, 32'd13821, -32'd2082, -32'd8121},
{-32'd9377, -32'd19785, -32'd1396, -32'd2755},
{32'd5125, -32'd12414, 32'd13752, 32'd2517},
{-32'd5787, -32'd3879, 32'd5566, 32'd1462},
{-32'd5437, 32'd7313, 32'd4054, 32'd5536},
{-32'd3424, -32'd5756, 32'd4326, 32'd6627},
{-32'd5630, -32'd2387, 32'd4387, 32'd2864},
{-32'd10032, 32'd7148, 32'd6829, -32'd2264},
{-32'd4943, 32'd7115, -32'd3032, -32'd2182},
{-32'd6078, -32'd3670, -32'd10583, -32'd9219},
{32'd5442, -32'd594, 32'd9947, 32'd3330},
{-32'd3318, 32'd2415, -32'd4600, -32'd91},
{32'd9415, 32'd10063, -32'd3372, -32'd6223},
{-32'd3210, 32'd239, 32'd2544, -32'd217},
{-32'd630, -32'd9274, -32'd9319, -32'd575},
{-32'd7492, 32'd9927, 32'd6440, -32'd5082},
{-32'd10705, -32'd1866, 32'd1807, 32'd14809},
{32'd10926, -32'd12862, -32'd18710, -32'd4102},
{32'd3626, 32'd9478, -32'd651, -32'd2899},
{-32'd2406, -32'd3181, 32'd9569, 32'd928},
{-32'd8765, -32'd2529, 32'd6092, 32'd3677},
{-32'd363, 32'd14678, 32'd2292, -32'd2131},
{32'd2734, 32'd13857, 32'd7372, 32'd10223},
{-32'd711, -32'd1428, -32'd4190, 32'd2350},
{32'd5159, -32'd111, 32'd1955, -32'd16166},
{-32'd8467, -32'd2595, 32'd612, 32'd3764},
{-32'd156, 32'd11278, 32'd7909, -32'd3467},
{32'd952, -32'd7369, -32'd7035, 32'd10654},
{32'd8394, 32'd4087, -32'd1104, 32'd2231},
{32'd3672, -32'd6929, -32'd12141, -32'd4354},
{32'd4957, -32'd445, -32'd1497, -32'd144},
{32'd7423, -32'd14822, -32'd13343, 32'd1099},
{-32'd4066, -32'd4934, 32'd5966, 32'd5774},
{32'd12990, 32'd3210, 32'd3824, 32'd8540},
{-32'd3918, -32'd4918, -32'd11130, -32'd5299},
{-32'd12707, 32'd5407, -32'd5903, 32'd4395},
{-32'd2184, 32'd16311, 32'd8870, -32'd5633},
{-32'd2077, 32'd2393, -32'd1193, 32'd7307},
{32'd9283, 32'd12220, -32'd96, 32'd653},
{-32'd6532, 32'd6834, 32'd218, 32'd1476},
{-32'd2780, -32'd4556, -32'd10432, -32'd3293},
{-32'd2316, 32'd989, 32'd8728, 32'd13038},
{-32'd9168, 32'd5640, -32'd10686, -32'd5570},
{-32'd3481, 32'd2542, -32'd4875, -32'd8895},
{32'd901, 32'd10406, -32'd2343, -32'd4773},
{-32'd467, -32'd871, 32'd5588, 32'd7180},
{32'd2120, 32'd1233, 32'd5243, -32'd11770},
{32'd9862, 32'd848, -32'd495, 32'd3418},
{32'd16000, 32'd3837, -32'd3505, -32'd6932},
{32'd3880, 32'd1901, -32'd2403, 32'd157},
{32'd3371, 32'd159, -32'd3495, -32'd1991},
{32'd6138, 32'd13793, 32'd6147, -32'd11310},
{32'd1897, 32'd3515, 32'd5094, 32'd8416},
{-32'd1082, 32'd1601, 32'd6644, 32'd5250},
{-32'd6876, 32'd11001, 32'd3790, -32'd695},
{32'd8318, -32'd4993, -32'd15994, 32'd244},
{32'd10464, 32'd12139, -32'd3181, 32'd1446},
{-32'd1840, -32'd9935, -32'd6810, 32'd4349},
{32'd11511, 32'd5940, -32'd4616, 32'd6414},
{-32'd9767, 32'd3181, -32'd2290, -32'd1558},
{32'd2268, -32'd10816, -32'd13319, -32'd5859},
{-32'd6682, 32'd7021, 32'd10213, 32'd1048},
{-32'd4401, 32'd6169, 32'd711, 32'd47},
{-32'd16222, 32'd2294, 32'd3956, -32'd7385},
{32'd4795, -32'd5274, 32'd3397, 32'd2780},
{32'd3692, 32'd2038, -32'd10640, 32'd1320},
{-32'd4191, -32'd5801, -32'd6899, -32'd9764},
{32'd2145, 32'd12520, -32'd5982, -32'd10643},
{-32'd2161, -32'd452, -32'd3688, -32'd3951},
{32'd1512, 32'd8264, 32'd1850, 32'd11974},
{-32'd4007, 32'd4619, 32'd7045, -32'd5043},
{-32'd1060, 32'd9392, -32'd5708, -32'd14453},
{32'd7532, -32'd13692, -32'd2162, 32'd1575},
{-32'd4605, -32'd1948, -32'd14218, 32'd15183}
},
{{-32'd2408, 32'd14864, 32'd3130, -32'd701},
{32'd2930, -32'd14688, -32'd8166, -32'd5135},
{32'd3888, -32'd11011, -32'd4641, -32'd1556},
{32'd2699, -32'd4067, 32'd9515, 32'd9334},
{32'd9426, -32'd3707, 32'd5251, 32'd1173},
{-32'd3956, 32'd1084, -32'd2284, 32'd3142},
{32'd10981, -32'd1345, -32'd1985, -32'd5769},
{32'd2252, -32'd2499, -32'd14005, -32'd6703},
{-32'd19806, -32'd4567, 32'd3053, 32'd8942},
{32'd10074, 32'd5656, 32'd13211, 32'd10487},
{-32'd12291, -32'd9815, -32'd2726, -32'd2550},
{-32'd2032, 32'd344, 32'd3600, 32'd401},
{-32'd4513, -32'd7095, -32'd700, 32'd3030},
{-32'd13928, 32'd4898, 32'd3337, -32'd1947},
{32'd7055, -32'd2498, -32'd3932, -32'd4643},
{-32'd40, 32'd8463, -32'd298, -32'd1890},
{32'd1118, -32'd7872, -32'd3526, 32'd2059},
{-32'd199, 32'd7825, 32'd270, 32'd616},
{32'd7109, -32'd2175, 32'd431, -32'd4912},
{-32'd3409, 32'd2740, -32'd3495, -32'd4104},
{-32'd8434, 32'd2293, -32'd4217, 32'd9773},
{-32'd5817, -32'd7718, -32'd12284, 32'd1064},
{32'd7057, 32'd2530, 32'd2176, -32'd24},
{32'd3471, 32'd376, -32'd8470, -32'd1876},
{32'd11577, 32'd15323, 32'd4556, 32'd3154},
{32'd331, -32'd8925, -32'd10277, 32'd1347},
{32'd6738, -32'd118, -32'd2424, -32'd4242},
{32'd8102, -32'd2497, 32'd5572, 32'd2009},
{32'd265, 32'd5465, -32'd5892, 32'd1998},
{32'd8632, -32'd10479, -32'd1891, -32'd4107},
{-32'd5853, 32'd4587, -32'd3998, -32'd13126},
{-32'd8387, -32'd2035, -32'd5441, -32'd7627},
{-32'd1686, 32'd4206, 32'd13811, 32'd628},
{32'd8308, 32'd3119, 32'd1488, 32'd6355},
{32'd17217, 32'd3452, 32'd5067, 32'd3512},
{-32'd16315, -32'd7005, -32'd1651, 32'd5005},
{-32'd1539, -32'd4618, -32'd1207, -32'd859},
{-32'd10280, 32'd678, -32'd3018, -32'd1250},
{32'd3695, -32'd739, 32'd5140, -32'd887},
{-32'd1080, 32'd6132, 32'd91, -32'd5034},
{-32'd3440, -32'd982, -32'd949, -32'd4443},
{32'd2281, -32'd2369, 32'd5367, -32'd1475},
{-32'd3842, -32'd655, 32'd9601, 32'd2962},
{32'd9912, 32'd284, 32'd2626, -32'd2607},
{-32'd12395, -32'd1387, -32'd4162, -32'd6867},
{-32'd540, -32'd4286, 32'd6752, 32'd8152},
{32'd1888, -32'd5953, 32'd5405, -32'd4790},
{32'd3365, -32'd12397, -32'd2284, -32'd5098},
{32'd7231, 32'd11228, 32'd4287, -32'd3258},
{32'd8461, -32'd5016, -32'd75, -32'd2734},
{-32'd10018, -32'd7570, 32'd6875, -32'd3030},
{32'd12715, 32'd8453, -32'd2763, 32'd650},
{-32'd7579, 32'd5525, 32'd10023, -32'd2268},
{-32'd4596, -32'd8784, 32'd1550, -32'd2107},
{32'd9448, -32'd2537, 32'd2433, 32'd1725},
{-32'd3371, 32'd371, -32'd2377, -32'd5074},
{32'd11123, 32'd2217, 32'd1823, 32'd769},
{-32'd6753, 32'd706, -32'd9859, -32'd5613},
{-32'd988, 32'd2728, -32'd5147, -32'd6357},
{-32'd3896, 32'd9179, 32'd4147, -32'd6805},
{32'd4885, -32'd4788, 32'd1850, -32'd1480},
{-32'd1849, -32'd13426, -32'd1155, 32'd7740},
{-32'd19910, -32'd8006, -32'd7348, -32'd4871},
{32'd3795, 32'd458, -32'd2820, -32'd3047},
{32'd7275, 32'd2014, -32'd1098, -32'd5},
{32'd4455, 32'd649, 32'd6176, 32'd2385},
{32'd8013, 32'd5991, -32'd862, 32'd341},
{32'd17558, -32'd789, -32'd5178, -32'd2829},
{32'd592, -32'd2883, -32'd453, 32'd674},
{32'd3813, -32'd2735, -32'd11636, 32'd2088},
{-32'd3865, 32'd1528, 32'd40, -32'd5093},
{32'd4143, -32'd7295, -32'd724, 32'd589},
{32'd10720, 32'd15, -32'd1258, -32'd12791},
{32'd15965, -32'd2743, -32'd5287, -32'd305},
{32'd2711, 32'd143, -32'd3381, 32'd3704},
{-32'd2347, -32'd419, 32'd2821, -32'd3536},
{32'd1226, -32'd15488, -32'd2304, -32'd3889},
{-32'd139, 32'd8133, -32'd7300, 32'd414},
{32'd7021, -32'd1904, 32'd8917, 32'd6572},
{-32'd6888, -32'd2284, -32'd3194, -32'd4535},
{32'd5607, 32'd7544, 32'd6328, 32'd5615},
{32'd7854, 32'd4985, 32'd1554, 32'd2432},
{-32'd1626, -32'd7244, -32'd338, -32'd6153},
{-32'd2552, 32'd7413, -32'd3786, -32'd5396},
{-32'd7513, 32'd6795, 32'd4468, -32'd2170},
{32'd5118, 32'd4613, -32'd2384, 32'd414},
{-32'd2153, -32'd438, 32'd2281, 32'd1977},
{-32'd173, -32'd4844, -32'd5437, -32'd6309},
{32'd4232, 32'd1038, -32'd2321, 32'd4082},
{-32'd378, 32'd3151, -32'd4784, -32'd5324},
{32'd6661, 32'd5277, 32'd5754, 32'd1043},
{-32'd2007, -32'd3523, -32'd4155, -32'd1190},
{32'd7279, 32'd4720, 32'd1716, -32'd742},
{32'd5286, 32'd5576, -32'd1084, 32'd4257},
{-32'd8463, -32'd5284, -32'd1074, 32'd3358},
{-32'd1273, 32'd1942, 32'd3550, -32'd4885},
{32'd5637, -32'd402, 32'd4520, 32'd1548},
{-32'd12232, 32'd4535, -32'd4888, -32'd2490},
{-32'd1841, -32'd4702, -32'd2677, -32'd7418},
{32'd6831, 32'd2963, 32'd6057, 32'd6249},
{32'd226, -32'd2785, 32'd5555, 32'd307},
{-32'd5876, 32'd892, -32'd5730, -32'd1781},
{32'd4238, -32'd5306, -32'd2578, -32'd2137},
{32'd4762, -32'd515, 32'd3959, 32'd928},
{-32'd1860, 32'd8213, 32'd690, 32'd1941},
{32'd8250, -32'd7486, -32'd2863, 32'd3465},
{-32'd2737, -32'd3195, -32'd14204, -32'd3848},
{-32'd4163, -32'd83, 32'd1866, 32'd875},
{32'd3214, 32'd6625, 32'd7531, 32'd3946},
{-32'd12826, 32'd3985, 32'd5457, -32'd6520},
{32'd3867, -32'd1733, 32'd4758, -32'd3400},
{32'd2713, 32'd2604, 32'd6229, 32'd5411},
{32'd14192, 32'd4819, 32'd8228, 32'd450},
{32'd11315, 32'd17039, -32'd1758, -32'd1644},
{-32'd4824, -32'd7171, -32'd2476, -32'd3444},
{32'd2365, 32'd596, 32'd2667, -32'd4742},
{32'd12404, -32'd6403, -32'd6021, -32'd381},
{-32'd4460, -32'd2245, 32'd2568, -32'd4504},
{-32'd223, 32'd16155, -32'd3072, 32'd6195},
{-32'd1707, 32'd5740, 32'd9658, -32'd813},
{32'd3186, -32'd6014, 32'd5849, -32'd1395},
{-32'd9324, -32'd7591, 32'd7817, 32'd3575},
{32'd6710, -32'd255, 32'd13289, 32'd1246},
{32'd1673, -32'd4794, -32'd5877, 32'd7532},
{32'd1338, -32'd4961, -32'd5130, 32'd713},
{32'd5780, 32'd2780, -32'd1916, 32'd1040},
{-32'd7960, -32'd4075, 32'd4339, -32'd3446},
{32'd1274, -32'd12052, 32'd2551, -32'd634},
{-32'd4674, -32'd7861, -32'd7524, -32'd2600},
{-32'd8339, -32'd820, -32'd3706, -32'd7106},
{-32'd3303, 32'd12886, -32'd4562, 32'd411},
{-32'd1822, -32'd3539, -32'd8942, -32'd10662},
{-32'd11373, 32'd2488, -32'd4787, -32'd1916},
{32'd4739, 32'd106, 32'd7726, -32'd1366},
{32'd5394, -32'd6350, -32'd383, 32'd3455},
{-32'd9371, 32'd8938, 32'd10574, 32'd2927},
{-32'd6855, -32'd5897, 32'd3061, -32'd882},
{-32'd8187, 32'd3509, 32'd3056, -32'd696},
{32'd7567, 32'd3896, -32'd2086, 32'd3913},
{32'd30, -32'd6407, -32'd6942, -32'd1464},
{-32'd8176, 32'd11382, 32'd514, 32'd5078},
{-32'd8274, -32'd4716, -32'd2830, -32'd4670},
{32'd3870, -32'd2467, 32'd1983, 32'd4136},
{-32'd3977, -32'd13491, -32'd4523, -32'd12445},
{32'd6723, -32'd5355, 32'd13173, 32'd7300},
{32'd19979, 32'd7344, 32'd3764, 32'd3529},
{-32'd11623, 32'd46, 32'd1514, -32'd2666},
{-32'd10145, -32'd4105, -32'd3963, -32'd9326},
{-32'd656, 32'd1625, 32'd2146, 32'd9630},
{32'd4054, -32'd4443, -32'd7479, -32'd7339},
{-32'd2401, -32'd4344, -32'd5646, -32'd4058},
{32'd5294, 32'd1086, 32'd9628, 32'd3773},
{-32'd30277, -32'd3323, -32'd34, 32'd2913},
{32'd7299, -32'd4846, -32'd1270, -32'd6502},
{-32'd5392, -32'd4202, -32'd4099, -32'd9295},
{-32'd1901, -32'd5284, 32'd2886, 32'd9360},
{32'd9818, 32'd17080, 32'd1542, 32'd3632},
{32'd13045, -32'd2120, -32'd6843, 32'd2633},
{32'd15333, -32'd1228, 32'd479, 32'd1848},
{-32'd10004, 32'd4753, -32'd655, 32'd198},
{-32'd11498, -32'd18714, -32'd2058, 32'd3352},
{32'd620, 32'd4702, -32'd807, 32'd1788},
{-32'd16054, 32'd1131, 32'd1714, -32'd9083},
{32'd15085, -32'd4250, 32'd146, 32'd7015},
{-32'd5886, 32'd3537, 32'd2297, 32'd14030},
{-32'd110, -32'd4767, -32'd456, -32'd715},
{-32'd13430, -32'd1466, -32'd3475, 32'd4946},
{-32'd11291, -32'd2197, -32'd4374, -32'd4581},
{-32'd7031, -32'd1411, 32'd5620, 32'd3202},
{-32'd16979, -32'd205, -32'd8813, -32'd3774},
{-32'd4827, 32'd3377, -32'd15848, -32'd5204},
{32'd5371, 32'd6074, -32'd1051, -32'd2964},
{32'd13933, 32'd2371, 32'd8195, 32'd6379},
{-32'd1084, -32'd9068, 32'd1759, -32'd1865},
{32'd838, 32'd5831, 32'd1166, 32'd4944},
{-32'd5084, 32'd2382, 32'd1381, 32'd384},
{-32'd3125, -32'd4097, 32'd2878, 32'd5345},
{32'd11423, 32'd8475, 32'd7213, 32'd4615},
{-32'd1183, 32'd5327, -32'd8862, 32'd2737},
{32'd6737, -32'd8830, -32'd4836, -32'd5337},
{32'd8048, 32'd2469, -32'd1182, 32'd118},
{-32'd1991, -32'd7130, 32'd1000, -32'd3880},
{-32'd5021, -32'd4503, 32'd4218, -32'd2304},
{-32'd7638, -32'd9342, -32'd2795, 32'd1220},
{-32'd265, -32'd2274, 32'd926, 32'd7458},
{32'd7588, 32'd2245, 32'd297, -32'd5360},
{32'd10991, 32'd4810, 32'd2750, 32'd4270},
{32'd9546, -32'd1235, 32'd4035, -32'd1438},
{-32'd4450, -32'd9170, -32'd533, 32'd4010},
{32'd5530, -32'd7678, 32'd4136, 32'd2866},
{32'd10355, 32'd4511, -32'd4292, 32'd20},
{-32'd8171, -32'd1541, -32'd2353, -32'd3555},
{32'd3811, 32'd2680, -32'd5682, 32'd641},
{32'd1815, 32'd4799, 32'd7507, -32'd3370},
{32'd1708, 32'd2465, -32'd1298, 32'd2389},
{32'd2706, 32'd3616, -32'd435, -32'd11712},
{32'd5728, -32'd1159, -32'd2040, -32'd5734},
{-32'd7208, -32'd1750, 32'd4167, -32'd3242},
{-32'd535, -32'd8738, 32'd275, -32'd979},
{-32'd6115, -32'd1149, 32'd7354, 32'd2981},
{-32'd8942, -32'd3839, -32'd7719, -32'd5917},
{32'd2322, 32'd5321, -32'd4297, -32'd1772},
{32'd6544, -32'd2275, -32'd3075, 32'd192},
{32'd18601, -32'd6143, 32'd3375, 32'd5285},
{32'd4154, -32'd2046, -32'd927, -32'd1660},
{32'd2878, -32'd11408, 32'd5115, -32'd5018},
{32'd7281, -32'd6319, -32'd7983, 32'd4105},
{-32'd1484, -32'd415, 32'd1854, -32'd394},
{32'd1881, -32'd2681, 32'd2537, 32'd3718},
{-32'd6465, -32'd1282, 32'd1017, -32'd24},
{-32'd5782, -32'd8492, -32'd1381, -32'd8801},
{32'd7336, 32'd4826, 32'd1752, -32'd3414},
{-32'd5237, -32'd12847, -32'd5912, 32'd2306},
{-32'd12076, -32'd181, -32'd4458, 32'd10239},
{-32'd7255, 32'd133, 32'd2788, 32'd506},
{32'd7949, -32'd5159, -32'd1390, -32'd2150},
{32'd6419, 32'd6650, -32'd3753, -32'd2517},
{-32'd197, -32'd13103, -32'd11757, 32'd955},
{32'd2039, 32'd17606, -32'd6612, -32'd2169},
{32'd2051, -32'd4427, -32'd3922, 32'd1814},
{32'd12543, 32'd2979, 32'd5744, -32'd1325},
{32'd1388, -32'd2104, -32'd1961, 32'd691},
{32'd1429, -32'd3179, 32'd4698, -32'd3358},
{32'd4413, 32'd4913, 32'd2990, -32'd2442},
{-32'd11256, -32'd1886, -32'd2927, -32'd264},
{32'd8620, 32'd1575, -32'd976, -32'd593},
{32'd9902, -32'd6298, -32'd4700, 32'd6620},
{-32'd6359, -32'd10014, 32'd66, 32'd4476},
{32'd1299, 32'd11624, -32'd1277, 32'd8423},
{-32'd3064, 32'd1428, -32'd342, 32'd2575},
{32'd2661, 32'd1595, -32'd2573, 32'd7320},
{32'd3757, -32'd8186, 32'd3932, -32'd176},
{32'd2159, 32'd3509, 32'd1515, -32'd4907},
{-32'd3462, -32'd16504, 32'd1779, 32'd2082},
{32'd7493, 32'd1421, 32'd368, -32'd1698},
{32'd1580, -32'd15904, 32'd1752, -32'd7265},
{32'd2766, -32'd4973, 32'd0, 32'd4722},
{32'd6326, -32'd7839, 32'd1689, -32'd4879},
{-32'd4819, 32'd675, 32'd9311, 32'd2629},
{32'd2056, -32'd11510, -32'd3735, -32'd3977},
{-32'd1670, 32'd2511, -32'd3840, -32'd1329},
{32'd1678, -32'd6704, -32'd2747, 32'd6902},
{-32'd10130, -32'd21492, -32'd12731, -32'd12240},
{-32'd10914, 32'd6453, 32'd4086, 32'd8963},
{32'd6972, 32'd8716, 32'd12182, 32'd6855},
{32'd7351, 32'd742, 32'd769, -32'd4169},
{32'd5829, -32'd2047, -32'd2868, -32'd6897},
{32'd4030, 32'd4748, 32'd1228, -32'd7062},
{32'd3324, -32'd6546, -32'd12257, 32'd3617},
{-32'd12383, -32'd14651, -32'd5385, 32'd1791},
{32'd3202, -32'd1899, -32'd747, 32'd6100},
{32'd9802, -32'd2905, -32'd832, -32'd5077},
{32'd3019, 32'd9370, 32'd7022, -32'd354},
{-32'd78, 32'd2547, -32'd5974, 32'd1794},
{-32'd4392, -32'd9582, -32'd6841, -32'd6519},
{32'd9051, -32'd3416, -32'd1177, 32'd979},
{32'd13478, -32'd5193, -32'd3999, 32'd1289},
{-32'd3650, -32'd1380, 32'd2074, 32'd4095},
{-32'd986, -32'd11281, -32'd10625, 32'd3129},
{-32'd7729, 32'd12208, 32'd2949, -32'd5204},
{32'd10700, 32'd11885, -32'd1989, -32'd3772},
{32'd12766, 32'd12818, 32'd3549, 32'd7023},
{32'd10522, -32'd7184, -32'd6018, -32'd2868},
{32'd5194, -32'd4786, 32'd1555, -32'd1667},
{32'd6072, -32'd2028, -32'd6477, 32'd5137},
{-32'd4685, 32'd2349, 32'd6649, 32'd8803},
{-32'd1376, 32'd5443, 32'd3652, 32'd11732},
{-32'd6499, 32'd3377, 32'd4461, 32'd211},
{32'd7094, -32'd4728, -32'd3029, -32'd1752},
{32'd8097, -32'd4551, -32'd1210, 32'd4177},
{-32'd1067, 32'd7391, 32'd1047, 32'd1005},
{32'd8018, -32'd14250, -32'd272, 32'd6929},
{32'd4050, -32'd1262, 32'd3147, -32'd6165},
{-32'd6586, -32'd8688, -32'd3631, -32'd12002},
{-32'd3452, -32'd4539, 32'd90, 32'd1656},
{-32'd6876, -32'd1067, 32'd1309, -32'd11361},
{32'd6727, 32'd7581, 32'd13355, 32'd11256},
{-32'd9970, 32'd6864, 32'd2537, -32'd1812},
{-32'd4886, -32'd9361, -32'd11928, -32'd9936},
{32'd4415, 32'd12096, -32'd1005, -32'd3754},
{-32'd6695, 32'd5824, 32'd5032, 32'd5789},
{-32'd6647, 32'd7116, 32'd7214, -32'd2961},
{32'd884, 32'd7230, -32'd4702, 32'd6670},
{-32'd5177, -32'd2062, -32'd3696, -32'd3018},
{-32'd10662, 32'd4937, 32'd1782, -32'd884},
{-32'd3018, -32'd6876, -32'd8746, -32'd3678},
{-32'd479, 32'd11681, 32'd4254, 32'd254},
{-32'd4780, -32'd5591, 32'd172, -32'd3462},
{32'd3442, 32'd9293, 32'd2183, -32'd6240},
{32'd8413, -32'd5678, 32'd3061, -32'd3404},
{-32'd5159, -32'd15831, 32'd1538, 32'd4800},
{32'd5880, 32'd6678, 32'd9505, 32'd1693},
{-32'd5186, 32'd2897, -32'd1098, 32'd7962},
{32'd7279, -32'd7906, -32'd4911, 32'd4644},
{-32'd7332, -32'd889, 32'd3862, 32'd4782},
{-32'd2339, 32'd451, -32'd3284, -32'd7337},
{32'd8128, -32'd3654, 32'd900, 32'd3459},
{-32'd3008, 32'd1871, 32'd118, 32'd481},
{32'd1566, 32'd2961, 32'd14184, 32'd3506},
{-32'd1382, -32'd1982, -32'd688, -32'd3901}
},
{{32'd1790, 32'd23470, -32'd6252, -32'd8459},
{-32'd5683, 32'd4707, -32'd8701, 32'd1725},
{32'd7001, 32'd4299, 32'd2618, -32'd5314},
{32'd4740, 32'd1449, 32'd12206, 32'd7455},
{32'd162, 32'd2909, 32'd7970, 32'd2098},
{32'd5245, -32'd14049, 32'd831, 32'd681},
{-32'd2673, 32'd13314, 32'd5921, 32'd2901},
{32'd3296, 32'd2788, 32'd1814, -32'd3580},
{-32'd2969, -32'd7289, 32'd6807, 32'd9582},
{32'd4715, -32'd1516, 32'd14828, 32'd11816},
{-32'd9896, -32'd5690, 32'd1074, -32'd2445},
{32'd1927, 32'd8158, -32'd1558, -32'd6138},
{32'd6548, 32'd3015, 32'd2337, 32'd666},
{32'd5797, 32'd1483, 32'd3687, 32'd597},
{-32'd444, 32'd3012, -32'd6365, -32'd4875},
{-32'd4661, 32'd8221, -32'd11088, 32'd9167},
{32'd5551, 32'd10423, -32'd851, -32'd3524},
{32'd9454, 32'd17137, -32'd1884, -32'd12396},
{-32'd3499, 32'd1879, 32'd11964, 32'd8432},
{32'd2787, -32'd3850, 32'd135, 32'd2564},
{-32'd8086, 32'd5601, -32'd160, -32'd4738},
{-32'd8935, -32'd6846, -32'd899, -32'd5672},
{32'd8530, 32'd5736, -32'd1563, 32'd1358},
{-32'd14288, -32'd2711, -32'd2877, 32'd4270},
{32'd11800, -32'd10152, 32'd931, 32'd930},
{32'd7487, 32'd1856, -32'd3218, 32'd2021},
{32'd9395, 32'd8723, 32'd2672, 32'd6825},
{32'd150, 32'd7756, -32'd1521, 32'd808},
{-32'd18597, -32'd1502, 32'd4422, 32'd702},
{-32'd159, -32'd4694, -32'd4168, -32'd3160},
{32'd4151, 32'd1368, -32'd14553, 32'd1246},
{32'd2688, -32'd5279, -32'd6711, -32'd6846},
{-32'd929, 32'd7016, 32'd971, -32'd1996},
{-32'd947, -32'd357, -32'd6877, 32'd1750},
{32'd3908, -32'd1815, 32'd9518, 32'd12226},
{32'd1202, 32'd7801, 32'd8055, 32'd2745},
{-32'd9610, 32'd7397, -32'd5335, 32'd5936},
{-32'd9892, -32'd712, 32'd2896, 32'd2568},
{-32'd1163, 32'd5341, -32'd5628, -32'd1753},
{32'd693, 32'd8536, 32'd1896, 32'd5563},
{-32'd8938, 32'd2465, -32'd2786, -32'd7501},
{32'd5119, 32'd3582, 32'd5926, -32'd3942},
{32'd1240, 32'd6113, 32'd2000, 32'd3336},
{-32'd6920, 32'd458, -32'd5682, 32'd6275},
{-32'd482, -32'd1024, 32'd4034, 32'd3949},
{-32'd9389, -32'd11165, 32'd827, 32'd121},
{-32'd322, -32'd8669, 32'd9052, -32'd3549},
{32'd13859, -32'd7597, -32'd3564, -32'd1859},
{32'd9215, 32'd6853, 32'd3829, -32'd696},
{32'd7015, -32'd7202, 32'd240, -32'd2227},
{-32'd10629, 32'd153, -32'd2999, 32'd738},
{32'd3427, -32'd707, 32'd555, -32'd7977},
{32'd1217, 32'd4962, -32'd1741, -32'd5627},
{-32'd3131, 32'd112, 32'd6125, 32'd4346},
{-32'd11884, 32'd1242, -32'd6724, -32'd2782},
{32'd2918, 32'd1446, -32'd4825, -32'd7633},
{32'd13116, -32'd1033, 32'd174, 32'd1064},
{-32'd8629, 32'd713, -32'd12498, -32'd5119},
{-32'd9130, -32'd8028, -32'd2418, -32'd1917},
{32'd13409, 32'd8590, 32'd5947, 32'd2080},
{32'd4933, 32'd116, 32'd5628, 32'd2744},
{-32'd357, 32'd582, -32'd2007, -32'd3790},
{-32'd18576, 32'd393, -32'd2839, -32'd2928},
{32'd9795, -32'd15510, 32'd4677, -32'd3406},
{-32'd660, -32'd8609, -32'd2825, 32'd3865},
{32'd2616, 32'd4657, 32'd8713, 32'd758},
{32'd2833, -32'd5763, -32'd931, 32'd3057},
{-32'd1749, 32'd4654, -32'd1998, -32'd4836},
{32'd11987, -32'd3917, 32'd673, 32'd5174},
{32'd778, 32'd4897, 32'd1243, -32'd3122},
{-32'd10807, -32'd7297, -32'd6617, -32'd6472},
{-32'd12255, 32'd2616, -32'd3242, -32'd3679},
{-32'd1842, -32'd6965, -32'd8739, -32'd6497},
{32'd6126, 32'd7156, -32'd6820, 32'd1190},
{32'd1735, 32'd733, 32'd4070, -32'd1457},
{-32'd2437, 32'd12857, 32'd4462, 32'd301},
{32'd7272, -32'd22269, -32'd1578, -32'd8622},
{-32'd1767, -32'd3789, -32'd1000, 32'd6565},
{32'd9193, -32'd7301, -32'd2533, 32'd974},
{-32'd11162, 32'd2161, -32'd6152, -32'd5431},
{32'd6350, 32'd2259, -32'd3001, 32'd100},
{-32'd3320, 32'd11582, 32'd7448, 32'd11271},
{-32'd13927, -32'd9618, -32'd2618, -32'd66},
{-32'd6118, 32'd307, -32'd8979, -32'd7161},
{32'd91, 32'd3608, -32'd11402, -32'd3238},
{32'd6197, -32'd2709, -32'd3569, -32'd672},
{-32'd16714, 32'd7154, 32'd4583, 32'd4888},
{-32'd4279, -32'd3725, -32'd2311, 32'd254},
{-32'd2030, -32'd21391, 32'd2013, 32'd4928},
{32'd6421, 32'd1720, -32'd11584, -32'd7041},
{-32'd2982, 32'd9454, 32'd6021, 32'd6000},
{-32'd13802, 32'd1824, -32'd6574, -32'd6453},
{32'd3265, 32'd15319, 32'd2911, 32'd810},
{32'd3423, 32'd4816, 32'd6036, 32'd2239},
{-32'd4795, -32'd691, 32'd5299, 32'd5717},
{32'd3070, -32'd4879, -32'd558, -32'd1186},
{32'd983, 32'd1137, 32'd10041, 32'd247},
{32'd11774, 32'd2825, -32'd1315, -32'd5124},
{32'd5725, -32'd238, -32'd4703, -32'd3980},
{32'd4773, 32'd1786, 32'd8240, -32'd1979},
{-32'd9020, -32'd11399, -32'd2664, 32'd173},
{32'd3388, 32'd1948, -32'd6326, -32'd1770},
{-32'd12881, -32'd1832, 32'd3652, 32'd2454},
{-32'd3352, 32'd727, -32'd3473, -32'd6899},
{-32'd5273, -32'd4696, 32'd2513, 32'd8242},
{-32'd8336, -32'd2480, 32'd3720, 32'd3499},
{32'd9118, -32'd15630, 32'd4310, 32'd5093},
{32'd1244, -32'd9711, -32'd3246, 32'd3449},
{32'd3608, 32'd3999, 32'd1982, 32'd2353},
{32'd3190, -32'd4593, -32'd4770, -32'd1323},
{-32'd4281, 32'd2621, 32'd9316, 32'd7200},
{-32'd1650, -32'd9187, 32'd4554, -32'd2769},
{32'd14921, 32'd702, 32'd3323, -32'd2116},
{-32'd8824, 32'd17458, -32'd626, -32'd3755},
{-32'd7806, -32'd8431, 32'd573, 32'd7478},
{-32'd3194, -32'd7855, -32'd5081, -32'd3564},
{-32'd4262, -32'd13921, -32'd7812, 32'd3370},
{-32'd5431, -32'd14669, -32'd6465, -32'd5302},
{32'd1725, -32'd5276, -32'd3804, 32'd974},
{32'd6590, 32'd1137, 32'd3400, 32'd2859},
{32'd1002, 32'd16068, -32'd385, 32'd10993},
{-32'd3478, -32'd2881, 32'd8427, -32'd4373},
{-32'd1685, 32'd13970, 32'd3348, -32'd4183},
{32'd5963, 32'd39, 32'd4497, 32'd4433},
{32'd721, 32'd878, -32'd3023, -32'd3690},
{32'd974, -32'd1388, -32'd777, -32'd5418},
{32'd15153, -32'd5702, 32'd5104, 32'd8791},
{32'd902, 32'd4853, -32'd2404, 32'd3914},
{-32'd13570, -32'd4188, 32'd1056, -32'd4196},
{-32'd10697, -32'd2848, -32'd11053, -32'd2203},
{-32'd1857, -32'd5629, -32'd362, -32'd497},
{32'd4061, -32'd5463, -32'd1814, 32'd1154},
{-32'd4392, -32'd8573, -32'd7733, -32'd534},
{32'd7761, 32'd3647, 32'd6583, -32'd3367},
{32'd5407, 32'd4776, 32'd7392, 32'd514},
{-32'd3322, -32'd425, -32'd9991, 32'd3533},
{-32'd10802, 32'd993, 32'd5363, 32'd2715},
{-32'd792, 32'd9839, -32'd2568, -32'd3802},
{32'd8523, -32'd1076, -32'd2224, 32'd6725},
{-32'd7309, 32'd2162, -32'd9507, -32'd5151},
{32'd1435, 32'd8118, 32'd6708, 32'd1123},
{-32'd10067, 32'd1121, -32'd4629, -32'd861},
{-32'd5349, -32'd2135, 32'd1747, -32'd7042},
{32'd1820, -32'd7938, -32'd7841, -32'd4707},
{32'd2455, 32'd7090, 32'd10289, 32'd789},
{32'd1316, 32'd16764, -32'd4234, 32'd5665},
{-32'd6880, -32'd11207, -32'd13015, 32'd3404},
{-32'd6159, -32'd159, -32'd9504, -32'd4384},
{32'd4484, 32'd5340, -32'd2428, -32'd6024},
{32'd5377, 32'd1987, -32'd5423, 32'd563},
{-32'd13745, 32'd4649, -32'd12836, 32'd1758},
{-32'd472, 32'd6322, 32'd9167, -32'd2298},
{-32'd10318, 32'd6559, 32'd2118, -32'd3852},
{-32'd2342, -32'd1361, -32'd3509, 32'd154},
{32'd122, -32'd5444, -32'd872, -32'd1616},
{-32'd4574, -32'd3847, -32'd3705, -32'd1056},
{32'd5118, 32'd5764, 32'd5948, 32'd2394},
{32'd1046, -32'd9870, -32'd6584, -32'd3458},
{-32'd7272, -32'd6304, 32'd1788, 32'd1686},
{32'd4375, -32'd3687, -32'd1560, 32'd3808},
{32'd6623, -32'd4895, 32'd4512, 32'd2025},
{32'd4953, -32'd4109, -32'd4857, 32'd13597},
{-32'd2269, -32'd8849, 32'd3368, -32'd2114},
{32'd4048, 32'd4135, -32'd3087, 32'd941},
{32'd538, 32'd3291, -32'd1164, -32'd3047},
{32'd7644, -32'd1649, -32'd6320, -32'd6638},
{-32'd11588, -32'd2778, 32'd1228, -32'd2866},
{-32'd1945, -32'd5972, -32'd780, 32'd2101},
{32'd2206, -32'd11705, 32'd2711, -32'd8217},
{-32'd13046, -32'd2753, -32'd13896, -32'd6258},
{-32'd3580, -32'd1923, 32'd1788, -32'd15647},
{32'd9710, 32'd4598, -32'd944, 32'd3969},
{32'd6928, 32'd6402, 32'd8760, 32'd9668},
{32'd2012, 32'd5188, -32'd3710, 32'd2793},
{32'd5895, -32'd5584, 32'd6716, -32'd13474},
{-32'd7253, -32'd19451, 32'd440, 32'd349},
{32'd1860, -32'd3369, -32'd1108, -32'd3178},
{32'd13919, 32'd2882, -32'd5448, -32'd244},
{32'd3182, 32'd14465, 32'd5356, 32'd9442},
{-32'd4593, 32'd2078, -32'd4147, -32'd5854},
{32'd2553, 32'd7856, -32'd8686, 32'd3304},
{-32'd7299, -32'd4005, -32'd147, 32'd2001},
{32'd4256, -32'd2658, -32'd4956, -32'd6619},
{-32'd9082, 32'd11158, -32'd5485, 32'd9144},
{-32'd5711, -32'd7841, 32'd13528, 32'd6489},
{32'd2030, 32'd2499, -32'd1387, 32'd305},
{32'd6312, 32'd13246, 32'd7364, -32'd5507},
{32'd760, 32'd8485, 32'd11183, 32'd8218},
{32'd6199, -32'd5033, 32'd2116, 32'd9212},
{-32'd3222, 32'd406, -32'd4159, 32'd2523},
{32'd1970, 32'd9981, -32'd9819, -32'd562},
{-32'd4070, -32'd8225, -32'd7540, 32'd2701},
{32'd10775, -32'd17326, 32'd9758, 32'd661},
{32'd7060, 32'd3846, -32'd2545, 32'd393},
{32'd8324, 32'd7691, 32'd1709, 32'd3098},
{-32'd5362, 32'd10829, 32'd5246, 32'd2220},
{-32'd898, 32'd3536, -32'd5179, -32'd4687},
{-32'd8604, 32'd5257, -32'd9647, 32'd1103},
{32'd3986, 32'd334, -32'd2215, 32'd5410},
{32'd5454, -32'd4972, -32'd3648, 32'd5622},
{-32'd3873, -32'd378, -32'd6289, -32'd4704},
{32'd1849, 32'd4592, -32'd11333, -32'd4151},
{-32'd4110, -32'd4768, -32'd809, 32'd9676},
{-32'd2480, 32'd3866, 32'd1500, 32'd2283},
{32'd937, -32'd7419, -32'd1380, 32'd4612},
{-32'd3851, -32'd1795, 32'd652, -32'd3691},
{32'd2562, -32'd2650, 32'd7058, -32'd729},
{-32'd11742, -32'd13400, -32'd1469, 32'd2346},
{32'd4364, 32'd11588, -32'd4755, -32'd2211},
{32'd2426, 32'd1271, -32'd6380, 32'd5722},
{32'd4577, 32'd2447, 32'd3976, -32'd565},
{32'd2215, -32'd7348, 32'd786, 32'd4362},
{32'd696, 32'd4426, -32'd3598, -32'd1219},
{32'd3693, -32'd3252, 32'd8509, -32'd1033},
{-32'd4057, 32'd5311, -32'd8372, 32'd6186},
{-32'd10225, -32'd4729, -32'd6067, -32'd1115},
{32'd4037, 32'd4675, 32'd5315, -32'd6253},
{-32'd6267, -32'd1699, -32'd3840, -32'd3705},
{-32'd7578, 32'd7594, -32'd8788, -32'd1209},
{-32'd2497, 32'd1071, -32'd2601, -32'd2594},
{-32'd4149, -32'd2484, -32'd4263, -32'd5057},
{32'd365, 32'd11644, 32'd2393, 32'd8143},
{-32'd6530, -32'd4767, 32'd10, 32'd8381},
{-32'd231, -32'd7302, -32'd6948, -32'd50},
{-32'd4688, -32'd5148, -32'd11384, -32'd1405},
{32'd2370, -32'd303, 32'd956, -32'd850},
{-32'd2120, -32'd442, -32'd3330, 32'd6596},
{32'd3182, -32'd5529, 32'd187, 32'd6233},
{32'd7749, 32'd10581, 32'd7975, 32'd8544},
{32'd4052, 32'd1728, -32'd1551, -32'd5960},
{-32'd3673, -32'd4171, -32'd10403, -32'd7185},
{-32'd1826, -32'd5714, -32'd5982, -32'd8093},
{32'd2016, 32'd7396, -32'd8592, -32'd1055},
{-32'd2204, 32'd19094, 32'd925, 32'd3914},
{-32'd1302, 32'd11425, -32'd4896, -32'd3164},
{32'd3476, -32'd10277, 32'd5842, 32'd5583},
{-32'd6590, -32'd13682, 32'd9092, 32'd4366},
{-32'd11168, -32'd4811, 32'd706, -32'd5786},
{32'd1952, -32'd7335, -32'd1995, -32'd8311},
{-32'd8774, 32'd6249, -32'd4016, 32'd2065},
{32'd3260, 32'd11658, -32'd42, 32'd3766},
{32'd13880, 32'd8647, -32'd5264, -32'd2215},
{32'd1529, -32'd2047, -32'd12417, -32'd4868},
{-32'd12303, 32'd3269, 32'd1606, 32'd13220},
{-32'd1024, -32'd4574, 32'd10621, 32'd4027},
{32'd6571, -32'd11995, 32'd3477, -32'd1769},
{-32'd13429, 32'd4111, -32'd7664, 32'd1411},
{32'd11107, -32'd7256, 32'd7942, 32'd630},
{-32'd10616, -32'd8427, -32'd1333, -32'd6005},
{-32'd6292, 32'd4892, -32'd1366, 32'd1926},
{-32'd13122, -32'd16789, -32'd194, -32'd1767},
{32'd2613, -32'd4220, 32'd8697, 32'd6077},
{32'd373, -32'd4553, 32'd769, 32'd4866},
{-32'd6977, 32'd10069, 32'd1805, -32'd135},
{-32'd10382, -32'd8275, -32'd8473, -32'd4307},
{32'd10013, -32'd1647, -32'd1986, -32'd6458},
{-32'd1509, -32'd761, 32'd4579, 32'd1794},
{32'd3219, 32'd2473, -32'd341, 32'd6357},
{-32'd8552, -32'd10654, -32'd540, -32'd5440},
{32'd11765, 32'd6256, -32'd5082, -32'd3061},
{32'd3810, -32'd5025, 32'd6735, -32'd9949},
{-32'd3498, -32'd11451, 32'd3426, 32'd1282},
{32'd8841, -32'd2351, -32'd8801, 32'd186},
{32'd7249, 32'd1904, -32'd5145, 32'd3454},
{32'd1032, -32'd8713, -32'd875, -32'd1630},
{-32'd1306, 32'd16549, 32'd5196, -32'd2483},
{32'd41, 32'd158, -32'd2072, 32'd7279},
{32'd9025, 32'd1780, -32'd9192, 32'd5566},
{32'd10975, -32'd5204, -32'd630, 32'd4504},
{32'd3161, 32'd2704, 32'd1135, -32'd1090},
{-32'd4883, -32'd3829, 32'd645, -32'd2592},
{32'd8050, 32'd1028, 32'd1404, -32'd507},
{-32'd988, -32'd9120, -32'd7996, -32'd7287},
{32'd15, -32'd3230, 32'd2530, -32'd7129},
{-32'd2806, 32'd1160, -32'd1352, 32'd1374},
{32'd559, 32'd2113, -32'd4825, -32'd2638},
{32'd4519, 32'd1258, 32'd14952, 32'd8960},
{-32'd9781, 32'd5790, -32'd4887, 32'd1828},
{-32'd4352, -32'd5599, -32'd6106, -32'd5238},
{-32'd1432, -32'd11677, -32'd2542, -32'd8947},
{32'd11587, -32'd4835, 32'd8516, 32'd9083},
{-32'd5961, -32'd5804, 32'd5296, -32'd982},
{-32'd1143, -32'd4162, -32'd3881, 32'd3806},
{32'd468, -32'd11941, 32'd2644, -32'd612},
{-32'd1297, 32'd12913, -32'd6990, -32'd3803},
{-32'd7759, 32'd5312, -32'd10512, 32'd2192},
{-32'd2029, 32'd9658, 32'd3576, 32'd6278},
{-32'd2626, -32'd16036, -32'd5072, 32'd734},
{32'd614, 32'd6934, -32'd609, 32'd488},
{32'd288, -32'd1972, -32'd2182, -32'd3092},
{-32'd6115, -32'd121, 32'd4420, 32'd7280},
{32'd4164, 32'd9689, 32'd5126, -32'd2139},
{32'd8723, -32'd9299, 32'd3506, 32'd183},
{-32'd9812, 32'd5204, -32'd1167, 32'd8381},
{-32'd5254, 32'd1389, -32'd7361, -32'd2033},
{-32'd44, 32'd5801, -32'd12836, 32'd1727},
{32'd3068, -32'd6275, 32'd4847, 32'd2938},
{32'd2038, -32'd10054, 32'd16314, 32'd5635},
{32'd3478, 32'd2792, 32'd7736, 32'd8448},
{32'd1359, -32'd6358, 32'd4091, 32'd5021}
},
{{32'd422, 32'd6337, -32'd2685, -32'd3669},
{32'd2554, -32'd8919, 32'd3980, 32'd2372},
{32'd6202, -32'd9925, -32'd3841, 32'd3836},
{32'd19968, -32'd3796, -32'd5819, -32'd5061},
{-32'd2303, 32'd15886, -32'd3645, -32'd714},
{32'd8654, -32'd5098, 32'd7671, 32'd2673},
{-32'd737, 32'd6756, 32'd1857, -32'd11167},
{-32'd1888, 32'd11327, -32'd4691, -32'd84},
{32'd2812, -32'd6957, 32'd5163, 32'd2409},
{32'd7044, 32'd3220, 32'd8151, -32'd7817},
{32'd2780, -32'd6805, 32'd5889, -32'd115},
{32'd3723, 32'd3273, -32'd696, -32'd1574},
{-32'd1250, -32'd1958, 32'd3136, 32'd7670},
{-32'd2361, 32'd1914, 32'd2628, 32'd1195},
{-32'd2858, 32'd688, -32'd3466, 32'd12167},
{-32'd1828, 32'd428, 32'd9219, 32'd9429},
{32'd9017, 32'd13214, 32'd5546, -32'd5203},
{32'd4789, 32'd3753, -32'd3931, 32'd7722},
{-32'd6465, -32'd13972, -32'd6083, -32'd6788},
{32'd383, -32'd3859, -32'd2811, -32'd9684},
{32'd1024, -32'd6277, -32'd1911, -32'd1451},
{-32'd8966, -32'd8996, -32'd10562, 32'd4168},
{-32'd4068, 32'd2858, 32'd1108, -32'd9119},
{-32'd11850, -32'd3076, -32'd3149, 32'd7928},
{32'd6343, 32'd4072, -32'd1848, -32'd5471},
{-32'd44, 32'd8049, -32'd805, 32'd4386},
{32'd2705, -32'd338, -32'd1068, 32'd55},
{32'd5994, 32'd7999, 32'd549, 32'd545},
{32'd6647, -32'd12192, -32'd3643, 32'd2912},
{32'd2122, 32'd4557, -32'd36, -32'd8283},
{-32'd733, 32'd8709, 32'd2212, 32'd8554},
{-32'd243, -32'd3054, -32'd3370, 32'd5874},
{32'd2567, -32'd1543, -32'd5095, -32'd7691},
{-32'd3698, 32'd10850, 32'd8222, 32'd11974},
{32'd2112, 32'd7421, -32'd1599, -32'd5549},
{-32'd2533, -32'd354, -32'd861, 32'd14208},
{-32'd2455, 32'd5426, -32'd707, 32'd6913},
{32'd4928, 32'd1386, 32'd2856, 32'd3580},
{32'd65, 32'd3033, -32'd4703, -32'd14482},
{-32'd2097, 32'd4186, -32'd11230, -32'd2836},
{32'd20721, -32'd12489, 32'd1337, -32'd4546},
{32'd3463, 32'd799, -32'd3237, 32'd2878},
{-32'd9751, 32'd13308, -32'd2222, -32'd2452},
{-32'd2544, 32'd2298, 32'd9220, -32'd3316},
{-32'd19099, -32'd2299, 32'd4303, 32'd8958},
{32'd5263, -32'd3172, 32'd6741, 32'd457},
{-32'd4223, -32'd9811, 32'd1125, 32'd19266},
{-32'd3283, 32'd1326, 32'd4768, 32'd6693},
{-32'd15629, 32'd5177, 32'd4808, -32'd5826},
{32'd4305, 32'd4562, -32'd1379, -32'd1940},
{32'd15189, 32'd2636, -32'd7853, -32'd3907},
{32'd3795, 32'd7303, 32'd10536, 32'd5002},
{-32'd10874, -32'd5756, 32'd9356, -32'd1629},
{-32'd5214, -32'd1404, -32'd11696, -32'd3533},
{-32'd6699, 32'd9037, 32'd11002, 32'd3985},
{32'd9735, -32'd3098, -32'd383, -32'd855},
{32'd1973, -32'd1469, -32'd4731, -32'd6660},
{-32'd821, -32'd1634, -32'd4122, -32'd1960},
{-32'd10872, -32'd6607, -32'd5509, 32'd6377},
{32'd2875, -32'd6666, -32'd5230, -32'd13821},
{-32'd5505, -32'd14059, 32'd1196, -32'd2126},
{-32'd880, 32'd4322, -32'd7280, -32'd2731},
{32'd1396, -32'd7893, -32'd2261, 32'd1565},
{-32'd7595, -32'd2509, -32'd5489, 32'd4360},
{32'd1054, 32'd3986, 32'd5053, 32'd1903},
{-32'd3608, 32'd4220, -32'd5226, -32'd10836},
{32'd3193, 32'd14021, 32'd3789, -32'd4042},
{-32'd1931, -32'd249, 32'd14359, 32'd4650},
{32'd14728, -32'd6085, 32'd3788, 32'd2435},
{-32'd2544, 32'd13167, -32'd11005, 32'd1884},
{32'd1452, -32'd3512, 32'd4483, -32'd4774},
{32'd700, -32'd2989, -32'd1280, 32'd5216},
{32'd2560, 32'd1081, 32'd1055, 32'd2594},
{-32'd3819, -32'd14446, 32'd6893, -32'd9245},
{32'd7010, -32'd1829, -32'd2974, -32'd7182},
{32'd5490, 32'd9776, 32'd8187, -32'd9484},
{32'd1192, -32'd6311, -32'd4993, 32'd3098},
{-32'd2811, -32'd3779, -32'd1495, 32'd11340},
{-32'd2848, 32'd7177, 32'd4038, -32'd2622},
{-32'd638, 32'd6539, -32'd3546, 32'd12656},
{32'd4253, 32'd2092, 32'd1089, -32'd7809},
{32'd5653, -32'd6452, 32'd8300, -32'd11162},
{-32'd3666, -32'd14426, -32'd6428, -32'd989},
{32'd9514, 32'd730, 32'd6155, -32'd7434},
{32'd53, -32'd1201, 32'd2637, -32'd2259},
{32'd8805, -32'd9121, -32'd7032, -32'd8531},
{-32'd4454, 32'd7459, 32'd4404, 32'd753},
{-32'd15118, -32'd8853, -32'd15402, 32'd4041},
{32'd10889, -32'd15183, -32'd3480, 32'd9273},
{32'd2356, -32'd1357, 32'd1647, -32'd4184},
{32'd3252, 32'd2907, 32'd6508, -32'd9480},
{-32'd6176, -32'd11659, 32'd1058, -32'd8747},
{-32'd6689, 32'd7402, 32'd12488, 32'd4676},
{-32'd2853, 32'd492, 32'd7669, -32'd14342},
{-32'd9826, -32'd4578, -32'd1537, 32'd3752},
{32'd4056, 32'd19516, 32'd3473, -32'd13758},
{-32'd4268, 32'd16066, 32'd4396, -32'd4075},
{-32'd6911, 32'd15610, -32'd4253, 32'd4344},
{-32'd7147, -32'd13478, -32'd8912, -32'd8600},
{-32'd569, 32'd15335, 32'd777, 32'd4761},
{-32'd17506, -32'd18933, 32'd9484, 32'd2732},
{32'd329, -32'd4651, -32'd3493, -32'd6522},
{-32'd7441, 32'd4958, 32'd644, -32'd5497},
{32'd2099, -32'd2246, 32'd7131, 32'd4746},
{-32'd3533, -32'd2936, -32'd8723, -32'd8120},
{-32'd19031, -32'd6745, -32'd2052, -32'd974},
{-32'd882, -32'd3813, -32'd398, 32'd7706},
{32'd7114, 32'd5772, 32'd391, -32'd4875},
{-32'd5230, 32'd10689, 32'd7804, 32'd6013},
{-32'd6554, 32'd3914, -32'd1401, 32'd5657},
{32'd2281, -32'd4076, 32'd3743, 32'd3917},
{-32'd319, -32'd8937, -32'd3657, -32'd9453},
{-32'd2351, 32'd2122, 32'd5171, -32'd5123},
{32'd3403, 32'd3261, -32'd8547, -32'd2798},
{-32'd670, -32'd11468, -32'd3974, -32'd652},
{32'd68, -32'd8966, 32'd2157, -32'd8967},
{32'd5994, -32'd3952, 32'd3900, 32'd10789},
{32'd12756, 32'd8490, 32'd5723, 32'd2761},
{32'd13180, -32'd243, -32'd2082, -32'd2099},
{-32'd6593, 32'd8255, 32'd1597, 32'd3228},
{-32'd231, 32'd6108, -32'd4218, -32'd8570},
{-32'd5114, -32'd8820, -32'd2739, 32'd8478},
{32'd586, 32'd652, 32'd5547, 32'd1275},
{32'd9469, -32'd5489, 32'd4418, -32'd6611},
{-32'd13638, -32'd7263, -32'd9279, 32'd1195},
{32'd3084, 32'd2632, 32'd9499, -32'd1789},
{32'd4484, -32'd1228, 32'd628, 32'd4389},
{-32'd10606, -32'd7439, -32'd8966, -32'd6006},
{32'd10153, -32'd3073, 32'd3203, 32'd2697},
{-32'd3690, -32'd978, -32'd10000, -32'd106},
{32'd2814, -32'd256, -32'd3323, -32'd1395},
{-32'd701, -32'd904, 32'd7204, 32'd7455},
{-32'd17080, -32'd1072, -32'd1200, 32'd6347},
{-32'd6067, -32'd2691, -32'd5267, 32'd882},
{-32'd11745, 32'd8988, -32'd2489, 32'd6916},
{32'd6323, 32'd5395, -32'd2089, -32'd6108},
{32'd6367, -32'd698, -32'd11354, 32'd1637},
{32'd7707, 32'd1516, -32'd9384, 32'd13780},
{32'd14028, -32'd1375, -32'd15104, -32'd2794},
{32'd2044, -32'd9493, -32'd773, -32'd4699},
{-32'd8132, -32'd4658, -32'd446, 32'd290},
{-32'd8059, -32'd416, -32'd5564, 32'd9675},
{32'd1273, 32'd3636, -32'd295, 32'd730},
{32'd5051, -32'd3453, 32'd7901, -32'd11981},
{-32'd717, 32'd7370, -32'd6544, -32'd3683},
{32'd11561, 32'd5711, 32'd971, -32'd9236},
{-32'd4403, -32'd4895, 32'd10629, 32'd4036},
{32'd10994, -32'd2092, 32'd1209, 32'd6101},
{32'd2526, 32'd2633, 32'd2053, -32'd9821},
{-32'd1183, -32'd9293, 32'd1656, 32'd1302},
{-32'd2670, 32'd2751, -32'd3433, 32'd13983},
{-32'd6006, 32'd5001, -32'd1920, -32'd1365},
{-32'd7337, -32'd7365, -32'd2892, -32'd7714},
{32'd2650, 32'd8009, 32'd12847, 32'd7335},
{-32'd7042, -32'd5936, -32'd935, 32'd9435},
{-32'd9321, -32'd2079, 32'd561, -32'd6907},
{-32'd5577, -32'd4972, -32'd10897, -32'd751},
{-32'd3837, -32'd4021, -32'd7035, 32'd2274},
{-32'd13848, -32'd17299, 32'd435, 32'd1905},
{32'd2181, -32'd1814, 32'd2434, 32'd6563},
{-32'd5434, -32'd851, 32'd4774, 32'd1648},
{-32'd2162, 32'd9976, 32'd1983, -32'd2535},
{-32'd2860, 32'd7308, -32'd9279, 32'd9201},
{-32'd1109, 32'd15750, 32'd583, -32'd5528},
{-32'd4662, -32'd5375, -32'd5851, 32'd425},
{32'd10697, -32'd6865, 32'd4796, -32'd14047},
{-32'd10969, 32'd2648, 32'd8365, 32'd101},
{32'd769, -32'd7667, -32'd5102, 32'd2954},
{32'd7450, 32'd890, 32'd6059, 32'd3009},
{32'd7061, 32'd3382, 32'd2522, 32'd7343},
{32'd8536, 32'd1367, -32'd4249, 32'd7486},
{-32'd4592, 32'd2832, -32'd8771, -32'd29},
{-32'd1599, 32'd3576, 32'd914, -32'd5785},
{-32'd7218, -32'd762, -32'd240, 32'd4072},
{32'd1471, 32'd6884, -32'd6542, -32'd4443},
{32'd5642, 32'd10387, 32'd2836, 32'd8005},
{32'd12069, 32'd9017, 32'd4173, -32'd7623},
{32'd11027, -32'd7247, 32'd81, -32'd251},
{-32'd4622, 32'd135, -32'd1455, -32'd9021},
{32'd2175, 32'd5598, -32'd5380, 32'd300},
{32'd3989, -32'd8650, 32'd6747, 32'd7216},
{-32'd6418, 32'd506, 32'd11020, 32'd7574},
{-32'd1437, -32'd15338, 32'd7115, -32'd7707},
{-32'd1215, -32'd6943, -32'd9444, -32'd1641},
{-32'd7433, -32'd669, 32'd6011, 32'd10025},
{32'd6563, -32'd7448, 32'd5217, -32'd9515},
{32'd2548, 32'd3150, -32'd10865, -32'd1866},
{32'd4816, 32'd5741, 32'd8025, -32'd571},
{-32'd13834, -32'd14059, 32'd2417, -32'd4325},
{-32'd2160, -32'd2009, -32'd7148, 32'd3871},
{-32'd5301, 32'd1234, -32'd2150, 32'd398},
{-32'd4889, 32'd3121, 32'd5543, 32'd12486},
{-32'd181, 32'd8233, 32'd1495, 32'd403},
{-32'd11836, -32'd4940, -32'd9237, 32'd1572},
{32'd11508, 32'd3148, -32'd1035, -32'd2137},
{-32'd4398, 32'd4126, -32'd4696, 32'd2047},
{-32'd5088, 32'd12660, 32'd6337, 32'd6763},
{32'd7391, -32'd5736, -32'd1121, -32'd5148},
{32'd4533, -32'd3694, -32'd6860, 32'd2293},
{-32'd722, 32'd13946, 32'd7089, -32'd10765},
{-32'd3573, -32'd6724, -32'd469, 32'd6034},
{32'd1019, 32'd3777, 32'd1939, 32'd1899},
{32'd738, -32'd1048, -32'd4877, -32'd1412},
{32'd2330, -32'd3868, 32'd2432, -32'd4794},
{32'd1117, 32'd13779, -32'd4826, -32'd2687},
{32'd1034, 32'd9485, -32'd13758, -32'd7450},
{-32'd6738, -32'd2411, 32'd1026, 32'd2120},
{32'd1177, -32'd5571, 32'd1038, -32'd1728},
{32'd8388, 32'd8683, -32'd6519, 32'd5115},
{-32'd5564, 32'd3855, -32'd6202, -32'd2670},
{-32'd2214, -32'd3493, -32'd5365, 32'd9384},
{32'd11183, 32'd4966, 32'd9346, -32'd5489},
{32'd2069, -32'd4104, -32'd6448, 32'd7127},
{32'd6986, -32'd9370, -32'd6024, -32'd5845},
{-32'd2477, 32'd7586, 32'd8757, -32'd1541},
{-32'd2250, -32'd2597, -32'd3032, -32'd2647},
{32'd1842, 32'd6717, -32'd8069, -32'd7101},
{32'd11784, 32'd7008, -32'd4638, 32'd6419},
{32'd11034, 32'd8693, 32'd3044, -32'd2748},
{32'd4188, -32'd1496, -32'd14924, -32'd10239},
{32'd7457, -32'd9112, 32'd5613, -32'd2689},
{-32'd2611, 32'd4577, -32'd14810, -32'd2677},
{-32'd5249, -32'd8114, 32'd2130, -32'd9939},
{32'd21095, -32'd5608, 32'd10690, 32'd7516},
{-32'd5436, -32'd5268, -32'd992, 32'd1622},
{-32'd8554, -32'd11340, -32'd1729, -32'd1033},
{32'd1756, 32'd6798, 32'd8693, -32'd7573},
{-32'd1647, -32'd1700, -32'd132, -32'd2316},
{32'd4324, -32'd1919, -32'd15717, -32'd4342},
{32'd2646, 32'd3282, 32'd4038, 32'd6119},
{32'd2929, -32'd14013, -32'd11031, 32'd7587},
{32'd1019, 32'd5153, 32'd8651, -32'd8715},
{32'd4845, -32'd12622, -32'd2184, 32'd15023},
{-32'd2867, 32'd1225, 32'd3118, -32'd173},
{32'd1455, 32'd4965, 32'd164, -32'd145},
{-32'd10268, -32'd2361, 32'd2916, 32'd10338},
{32'd6171, -32'd1139, 32'd10552, -32'd1705},
{-32'd570, -32'd9129, -32'd751, 32'd10186},
{32'd8927, 32'd11457, 32'd3205, 32'd3813},
{32'd5412, -32'd3692, 32'd4248, 32'd2733},
{-32'd19322, -32'd10740, -32'd14468, -32'd10466},
{32'd4022, -32'd5586, -32'd6627, 32'd2106},
{32'd3370, 32'd2846, 32'd2305, 32'd8688},
{32'd7665, -32'd2436, 32'd9267, 32'd1764},
{32'd2033, 32'd2825, 32'd6329, -32'd5072},
{-32'd8501, 32'd1062, -32'd5616, 32'd3451},
{32'd4608, 32'd4593, -32'd6046, 32'd1613},
{-32'd1722, 32'd2044, 32'd2691, -32'd217},
{-32'd7180, -32'd2322, 32'd596, 32'd6874},
{32'd4277, -32'd1153, 32'd7035, -32'd8298},
{32'd677, -32'd12219, 32'd2306, 32'd2114},
{32'd2510, 32'd7226, 32'd7736, -32'd6633},
{32'd1679, 32'd13741, 32'd14430, -32'd7645},
{32'd753, -32'd1994, 32'd2053, -32'd3579},
{32'd1557, 32'd639, 32'd10199, -32'd8284},
{32'd9149, -32'd1963, -32'd873, 32'd9},
{32'd4394, 32'd246, 32'd7294, -32'd699},
{32'd13357, 32'd5737, 32'd8328, 32'd937},
{-32'd2437, -32'd10856, 32'd3190, 32'd6648},
{32'd14130, 32'd4063, -32'd4939, 32'd5138},
{32'd6641, -32'd3765, 32'd6003, -32'd4900},
{-32'd1212, 32'd5007, -32'd5710, 32'd4156},
{-32'd9312, 32'd1353, 32'd1515, -32'd11104},
{32'd1973, -32'd1620, -32'd4254, 32'd9352},
{32'd1954, 32'd5117, 32'd955, 32'd507},
{32'd238, -32'd12161, 32'd9345, -32'd10982},
{32'd4413, 32'd5426, -32'd455, 32'd12975},
{-32'd3618, -32'd2516, -32'd13159, 32'd2512},
{32'd11159, -32'd4457, 32'd1927, -32'd7382},
{-32'd2558, -32'd2923, -32'd3180, 32'd12744},
{32'd5724, -32'd361, -32'd9325, -32'd3553},
{32'd3974, 32'd6633, -32'd5867, -32'd1381},
{-32'd3045, -32'd793, -32'd7177, -32'd1943},
{32'd445, -32'd4634, 32'd2754, 32'd6818},
{32'd1302, -32'd5907, 32'd5296, -32'd7936},
{32'd520, -32'd3001, -32'd6717, 32'd7052},
{32'd3348, 32'd6112, 32'd5896, -32'd7586},
{32'd8012, 32'd8692, 32'd8960, 32'd5802},
{-32'd683, 32'd1184, 32'd3885, 32'd9041},
{-32'd682, 32'd4835, -32'd4477, 32'd6602},
{-32'd5851, 32'd5242, -32'd8483, -32'd5203},
{-32'd9144, -32'd8977, 32'd1186, -32'd3007},
{32'd238, -32'd6326, 32'd3497, -32'd3785},
{-32'd4287, -32'd12008, -32'd5536, 32'd6485},
{-32'd1419, 32'd7892, -32'd657, -32'd15400},
{32'd776, 32'd667, 32'd4507, 32'd2505},
{32'd616, 32'd668, -32'd2717, -32'd10943},
{32'd6238, 32'd6866, -32'd494, 32'd9628},
{-32'd5493, 32'd11190, -32'd7808, 32'd6346},
{-32'd4714, -32'd8936, -32'd2769, -32'd3075},
{-32'd7746, -32'd5763, -32'd8211, 32'd9181},
{32'd1422, -32'd51, 32'd13619, -32'd1180},
{-32'd3658, 32'd1662, 32'd3357, -32'd3725},
{-32'd4029, -32'd8685, 32'd7567, 32'd4155},
{-32'd322, -32'd5807, -32'd942, -32'd3330},
{32'd2812, 32'd12863, -32'd1586, 32'd450},
{-32'd8300, 32'd1393, -32'd159, 32'd3587},
{-32'd1838, 32'd4761, 32'd2187, -32'd4500},
{32'd5413, 32'd7158, 32'd2258, -32'd9163},
{-32'd5418, -32'd16979, 32'd9409, 32'd14116}
},
{{-32'd1926, -32'd3866, 32'd13227, 32'd6134},
{32'd728, -32'd2153, -32'd11407, -32'd7894},
{-32'd6431, -32'd1217, 32'd3447, -32'd596},
{32'd9080, -32'd4166, -32'd4614, 32'd7057},
{32'd6380, 32'd952, 32'd7974, 32'd5039},
{32'd4418, -32'd7206, -32'd6476, -32'd5869},
{32'd979, -32'd782, 32'd338, -32'd1959},
{32'd3283, -32'd4570, -32'd3154, -32'd2626},
{32'd3992, 32'd2361, 32'd3039, 32'd1736},
{32'd8002, 32'd5748, 32'd5060, 32'd10087},
{32'd7854, -32'd11422, 32'd7244, -32'd4974},
{32'd4686, 32'd3669, 32'd2370, 32'd1617},
{32'd6029, -32'd5679, 32'd5980, 32'd1807},
{-32'd6107, -32'd6108, -32'd5210, 32'd8870},
{-32'd9487, -32'd22215, 32'd1148, 32'd908},
{-32'd3014, 32'd7828, 32'd2933, 32'd8905},
{32'd5934, 32'd5578, 32'd9683, -32'd3239},
{32'd2732, 32'd9081, -32'd5469, 32'd3601},
{32'd3521, -32'd6584, 32'd5984, 32'd8095},
{32'd1320, -32'd4976, 32'd4704, 32'd11652},
{-32'd5534, -32'd2841, -32'd3857, 32'd2908},
{-32'd3625, -32'd4588, -32'd4003, 32'd1455},
{32'd7935, 32'd1487, -32'd5104, -32'd6576},
{-32'd11297, -32'd38, -32'd2017, -32'd1524},
{32'd7887, 32'd4135, -32'd2740, -32'd6984},
{-32'd8626, 32'd13457, 32'd1969, 32'd414},
{-32'd5207, -32'd1915, -32'd14984, -32'd1169},
{32'd9141, 32'd474, -32'd89, 32'd2583},
{-32'd1526, 32'd1239, 32'd5140, 32'd4250},
{-32'd4745, 32'd2788, 32'd4520, 32'd4777},
{-32'd4064, -32'd8353, 32'd10572, -32'd659},
{-32'd7990, -32'd5611, -32'd309, -32'd1793},
{32'd8761, 32'd1880, 32'd6937, 32'd2710},
{-32'd6860, -32'd171, 32'd8853, 32'd1102},
{32'd11480, 32'd6041, -32'd6, 32'd4411},
{-32'd5096, -32'd1855, 32'd823, -32'd2149},
{-32'd2921, 32'd10119, 32'd5198, -32'd1700},
{-32'd328, 32'd2760, 32'd6189, 32'd7681},
{32'd5591, -32'd8012, 32'd2496, -32'd1494},
{-32'd1374, -32'd9932, 32'd3314, -32'd4684},
{32'd1780, -32'd1931, -32'd2168, -32'd8459},
{-32'd272, 32'd4111, 32'd8467, 32'd28},
{32'd3348, -32'd4021, -32'd958, 32'd3447},
{-32'd5117, -32'd10631, 32'd5515, 32'd3498},
{-32'd7125, 32'd1464, 32'd1111, 32'd7534},
{32'd6054, -32'd1226, -32'd3466, 32'd11178},
{-32'd4957, -32'd9185, -32'd1836, -32'd612},
{-32'd2674, 32'd3795, 32'd2402, 32'd3269},
{-32'd1357, 32'd3639, -32'd382, -32'd1749},
{-32'd412, -32'd4019, -32'd2913, -32'd1274},
{-32'd2732, 32'd4789, 32'd854, 32'd8256},
{-32'd1809, 32'd4542, -32'd725, -32'd1725},
{-32'd7009, -32'd4373, -32'd5146, 32'd3275},
{-32'd1115, -32'd1640, 32'd10169, -32'd5665},
{32'd13624, 32'd6607, 32'd703, 32'd1900},
{32'd3595, -32'd7686, -32'd6957, -32'd2283},
{32'd4971, 32'd5614, -32'd476, -32'd3337},
{-32'd10345, -32'd11159, 32'd6470, -32'd4416},
{-32'd14810, -32'd12096, -32'd8129, -32'd6685},
{-32'd4899, -32'd333, -32'd6492, -32'd4695},
{-32'd9145, -32'd3748, 32'd1059, 32'd8814},
{-32'd3329, -32'd4189, 32'd1824, 32'd3524},
{-32'd12857, -32'd12776, -32'd737, 32'd508},
{-32'd2912, 32'd4085, -32'd1000, -32'd2205},
{32'd7395, 32'd2943, 32'd7319, -32'd4187},
{32'd7829, 32'd5388, 32'd3217, -32'd170},
{-32'd2862, -32'd8163, -32'd3519, -32'd625},
{32'd3022, 32'd3462, -32'd2357, -32'd437},
{32'd12089, -32'd1406, 32'd3108, -32'd2105},
{-32'd5864, 32'd3599, -32'd5209, -32'd6751},
{32'd3485, -32'd11196, -32'd1912, 32'd5510},
{32'd2762, 32'd2168, 32'd1151, -32'd1687},
{-32'd11995, -32'd2610, -32'd5364, -32'd4974},
{32'd4880, -32'd2896, 32'd2738, -32'd2100},
{32'd5137, 32'd3115, 32'd3378, -32'd1422},
{32'd1439, 32'd1596, -32'd1202, 32'd7127},
{-32'd13323, -32'd6032, 32'd456, -32'd2514},
{32'd249, -32'd5629, -32'd4160, 32'd321},
{32'd14334, 32'd1476, 32'd459, 32'd1139},
{-32'd4826, 32'd3906, -32'd4912, -32'd2090},
{32'd8753, 32'd6636, 32'd5081, 32'd3198},
{32'd244, -32'd533, 32'd8743, 32'd2285},
{32'd3310, -32'd15315, -32'd6143, -32'd4956},
{32'd10292, -32'd4050, 32'd608, 32'd367},
{-32'd6664, -32'd1428, -32'd774, 32'd5358},
{-32'd1645, 32'd7970, 32'd8157, 32'd908},
{32'd4013, 32'd5579, 32'd897, 32'd9989},
{-32'd6128, -32'd3442, 32'd5158, -32'd7047},
{-32'd838, -32'd5605, 32'd753, 32'd4089},
{-32'd2648, -32'd3728, -32'd5375, -32'd7979},
{32'd2721, -32'd1765, 32'd691, 32'd6634},
{-32'd1536, 32'd1145, -32'd2671, -32'd3628},
{32'd14722, 32'd7740, 32'd9754, 32'd7451},
{32'd4824, 32'd8748, 32'd120, 32'd3793},
{-32'd3637, 32'd1787, -32'd4792, -32'd3772},
{-32'd3579, 32'd1085, -32'd2957, -32'd5745},
{32'd5260, -32'd3278, 32'd7830, 32'd7078},
{-32'd5669, 32'd9547, 32'd44, -32'd1026},
{32'd311, 32'd7702, -32'd2942, -32'd5576},
{-32'd988, -32'd2788, 32'd1518, 32'd10706},
{-32'd10002, 32'd1305, 32'd2832, -32'd5058},
{-32'd1239, -32'd2034, 32'd94, -32'd3068},
{-32'd3079, -32'd661, 32'd4426, -32'd10326},
{32'd8757, 32'd2374, -32'd1355, -32'd1332},
{32'd8059, 32'd2891, 32'd3217, -32'd5590},
{-32'd11355, 32'd3766, -32'd9725, 32'd1257},
{-32'd3549, -32'd529, -32'd1624, -32'd6007},
{-32'd2772, -32'd2954, -32'd3609, 32'd2612},
{32'd4765, -32'd6541, 32'd72, 32'd1251},
{-32'd9214, 32'd871, 32'd5046, 32'd4210},
{32'd586, 32'd1279, -32'd11527, -32'd6162},
{-32'd191, 32'd1688, 32'd346, -32'd7502},
{-32'd2534, 32'd4768, 32'd6204, -32'd120},
{-32'd2417, 32'd48, -32'd7000, 32'd2862},
{32'd1580, -32'd7318, 32'd395, 32'd371},
{32'd4757, -32'd5956, -32'd17551, 32'd131},
{32'd5430, 32'd6019, 32'd2749, 32'd720},
{32'd14184, 32'd2672, -32'd3692, 32'd4690},
{-32'd5240, -32'd8187, 32'd2793, 32'd2859},
{32'd4847, 32'd13880, 32'd2931, 32'd1971},
{32'd8953, 32'd1112, -32'd2633, 32'd415},
{32'd2356, 32'd2608, 32'd7100, -32'd1854},
{32'd7125, -32'd1640, 32'd5559, 32'd6975},
{32'd4930, -32'd3339, -32'd6116, -32'd7389},
{-32'd5699, -32'd8180, 32'd4765, 32'd849},
{32'd2538, 32'd3396, -32'd4139, 32'd4717},
{-32'd1258, -32'd2005, -32'd7837, -32'd8134},
{-32'd5787, -32'd1980, 32'd1941, 32'd1768},
{-32'd217, 32'd2411, -32'd7365, -32'd9554},
{-32'd7556, 32'd4713, 32'd3260, 32'd4977},
{32'd10307, 32'd1184, 32'd7860, 32'd7390},
{-32'd4649, -32'd7789, 32'd2728, 32'd1394},
{-32'd7536, -32'd1111, 32'd1391, -32'd4728},
{32'd6594, 32'd6382, -32'd401, -32'd2179},
{32'd7571, -32'd6166, 32'd721, -32'd5307},
{-32'd5000, 32'd2578, 32'd5859, -32'd7090},
{32'd7601, 32'd3473, 32'd12745, -32'd631},
{-32'd16068, 32'd1213, 32'd1057, -32'd5984},
{32'd5773, 32'd9250, -32'd8570, 32'd398},
{-32'd6752, 32'd482, -32'd10364, -32'd5010},
{32'd552, 32'd6336, 32'd10173, 32'd5519},
{-32'd21, -32'd3750, -32'd1775, -32'd5464},
{32'd147, -32'd2072, -32'd200, 32'd937},
{32'd2268, -32'd6143, -32'd173, 32'd1005},
{32'd3863, 32'd9046, 32'd5365, 32'd1760},
{32'd2292, -32'd1385, 32'd6404, -32'd1577},
{32'd1280, 32'd702, 32'd1320, 32'd431},
{-32'd2659, -32'd8906, 32'd9805, -32'd5867},
{-32'd11043, -32'd2930, -32'd8523, 32'd2429},
{-32'd9150, -32'd12863, -32'd6185, -32'd1561},
{-32'd4201, -32'd1986, 32'd2947, -32'd340},
{32'd7481, -32'd3385, 32'd8547, 32'd1713},
{-32'd1796, 32'd1741, -32'd4655, -32'd46},
{-32'd7820, 32'd4084, -32'd5814, -32'd695},
{-32'd6760, -32'd4524, -32'd3073, -32'd5941},
{32'd11207, 32'd4583, -32'd1715, -32'd3428},
{32'd8403, 32'd1053, 32'd2316, -32'd316},
{-32'd2952, 32'd10223, -32'd2396, -32'd5946},
{-32'd10538, -32'd636, -32'd6387, -32'd1813},
{-32'd3968, -32'd7203, 32'd3839, 32'd5513},
{32'd785, -32'd2326, 32'd1111, -32'd2591},
{32'd18869, -32'd5186, 32'd13792, -32'd241},
{-32'd4927, -32'd6714, -32'd9813, -32'd1177},
{32'd3899, 32'd2212, -32'd909, -32'd6541},
{-32'd766, 32'd7297, -32'd6033, 32'd1653},
{-32'd11168, -32'd8267, -32'd7156, -32'd3371},
{32'd1855, -32'd1109, 32'd2405, 32'd496},
{-32'd4092, -32'd10551, -32'd2828, 32'd904},
{-32'd9578, -32'd1039, 32'd5331, 32'd5161},
{-32'd6857, 32'd7904, -32'd5055, -32'd2763},
{-32'd11062, -32'd8263, -32'd9424, -32'd9154},
{-32'd3181, 32'd4206, -32'd6326, -32'd586},
{32'd11722, 32'd9363, 32'd3889, 32'd4385},
{-32'd133, 32'd6192, 32'd3323, -32'd4021},
{-32'd2954, -32'd6706, -32'd25, -32'd5696},
{-32'd2313, -32'd2566, 32'd5972, 32'd4556},
{-32'd1382, 32'd6867, 32'd2241, 32'd3426},
{-32'd7183, 32'd3476, -32'd179, -32'd2994},
{32'd3652, 32'd1513, 32'd2235, -32'd1730},
{-32'd4749, -32'd12889, 32'd1087, -32'd1069},
{-32'd8846, 32'd4121, 32'd10183, -32'd767},
{-32'd5498, -32'd9678, 32'd3363, 32'd5419},
{32'd2825, -32'd9632, -32'd7805, -32'd3074},
{32'd3282, 32'd865, 32'd9756, 32'd5622},
{-32'd2704, 32'd6127, 32'd3678, -32'd2946},
{32'd2608, 32'd3006, -32'd6630, -32'd1402},
{-32'd6332, -32'd3631, -32'd6692, 32'd4259},
{32'd6198, -32'd4159, 32'd3248, -32'd2090},
{32'd1572, -32'd2069, 32'd2170, -32'd7597},
{32'd1843, -32'd7166, 32'd2556, 32'd6823},
{-32'd2041, -32'd2841, 32'd5884, 32'd3107},
{-32'd6975, -32'd13983, -32'd218, -32'd5246},
{-32'd6409, -32'd1645, -32'd6565, -32'd9108},
{-32'd2146, 32'd6852, -32'd170, -32'd4775},
{32'd10927, 32'd9086, -32'd9963, 32'd1273},
{-32'd2924, -32'd1157, -32'd1672, 32'd2076},
{-32'd7378, 32'd436, -32'd5224, 32'd1501},
{32'd4840, 32'd6252, -32'd3354, 32'd1264},
{32'd2567, -32'd3924, -32'd813, 32'd413},
{-32'd224, -32'd943, -32'd2585, 32'd114},
{-32'd7015, -32'd10941, 32'd2496, -32'd3180},
{32'd4167, -32'd3084, 32'd1502, 32'd100},
{32'd2643, -32'd1385, 32'd3348, 32'd5315},
{32'd5378, -32'd3557, -32'd2611, 32'd2332},
{32'd1106, 32'd816, 32'd1413, -32'd4413},
{32'd5746, 32'd10033, -32'd2710, 32'd3843},
{32'd13335, -32'd3962, -32'd1614, 32'd4494},
{-32'd5624, 32'd5468, 32'd3684, -32'd6613},
{-32'd7073, -32'd60, -32'd6237, -32'd6310},
{32'd3201, -32'd1860, 32'd4048, 32'd6305},
{-32'd5879, 32'd6002, -32'd4524, -32'd9719},
{-32'd4279, 32'd6175, 32'd5221, 32'd4071},
{32'd628, -32'd1949, -32'd2472, -32'd1018},
{32'd3452, 32'd3361, -32'd2641, -32'd10315},
{-32'd846, -32'd5753, -32'd4056, 32'd6232},
{32'd2006, 32'd4070, 32'd1160, -32'd573},
{-32'd5343, -32'd2009, -32'd3113, 32'd349},
{32'd13323, -32'd5247, -32'd4580, -32'd1688},
{-32'd2228, 32'd4678, 32'd4055, 32'd3868},
{-32'd1202, -32'd5791, -32'd3076, -32'd2851},
{-32'd5633, -32'd6958, 32'd4937, 32'd2496},
{-32'd1716, 32'd5317, 32'd3260, -32'd3242},
{32'd5584, 32'd3202, 32'd1856, 32'd2341},
{-32'd11711, 32'd11797, -32'd7338, -32'd5442},
{32'd3506, -32'd2729, -32'd5861, -32'd1327},
{-32'd2078, 32'd15308, -32'd14478, 32'd1092},
{32'd4209, -32'd6364, 32'd5352, 32'd1038},
{32'd7029, 32'd2336, -32'd5388, -32'd1753},
{32'd5032, 32'd1423, 32'd3651, -32'd2597},
{32'd8592, -32'd3936, 32'd123, 32'd2155},
{-32'd8138, -32'd6127, -32'd8178, -32'd4325},
{-32'd7883, -32'd2975, 32'd2277, 32'd4896},
{-32'd6180, 32'd1992, -32'd57, -32'd1780},
{-32'd1162, -32'd1055, -32'd2972, 32'd6320},
{-32'd3181, -32'd2432, 32'd603, 32'd6631},
{32'd3869, -32'd1251, -32'd9771, -32'd1147},
{32'd4198, -32'd6264, -32'd3818, -32'd7104},
{-32'd351, -32'd2108, -32'd9247, 32'd1818},
{32'd5590, -32'd5614, 32'd4444, 32'd2462},
{-32'd9365, 32'd7790, -32'd895, -32'd489},
{32'd900, 32'd235, -32'd1946, -32'd82},
{-32'd5512, 32'd15140, -32'd9050, 32'd1904},
{-32'd5025, -32'd8792, -32'd4574, -32'd4698},
{32'd3665, 32'd264, -32'd1714, 32'd1628},
{32'd10794, 32'd4261, 32'd5524, 32'd7155},
{32'd1344, -32'd984, 32'd5913, -32'd2978},
{-32'd1879, -32'd6986, -32'd2367, -32'd3555},
{32'd9079, -32'd4588, -32'd10148, 32'd4128},
{32'd5216, 32'd7975, -32'd1808, -32'd2498},
{32'd312, -32'd5826, -32'd11634, 32'd866},
{-32'd11583, 32'd4945, 32'd5274, 32'd1479},
{-32'd406, 32'd5914, 32'd7527, 32'd2540},
{-32'd2600, 32'd10489, 32'd2713, 32'd14772},
{32'd12377, -32'd8099, 32'd72, -32'd2993},
{32'd4584, -32'd6139, 32'd3264, 32'd3390},
{-32'd9408, 32'd11227, 32'd4759, -32'd158},
{32'd3343, 32'd6280, -32'd3033, -32'd1707},
{32'd2058, 32'd15650, 32'd4525, 32'd4499},
{32'd1203, -32'd5392, 32'd1790, -32'd9192},
{32'd6781, 32'd7400, -32'd5851, 32'd4779},
{-32'd4419, 32'd587, -32'd5297, 32'd589},
{-32'd4601, -32'd5588, -32'd3778, -32'd3236},
{32'd854, 32'd1843, 32'd2412, 32'd588},
{-32'd4321, 32'd9849, -32'd7606, -32'd5074},
{32'd6055, 32'd15908, 32'd2361, -32'd1980},
{-32'd6861, 32'd1758, 32'd912, 32'd2843},
{32'd9105, -32'd1448, -32'd5891, -32'd2492},
{-32'd13338, -32'd182, -32'd366, -32'd8},
{-32'd13464, -32'd2658, -32'd5329, -32'd8235},
{-32'd3471, -32'd6627, -32'd2003, -32'd4229},
{32'd8856, -32'd5487, 32'd2253, -32'd1195},
{32'd11099, 32'd8501, -32'd2470, -32'd12919},
{32'd1870, -32'd5129, 32'd8162, -32'd3158},
{32'd5013, -32'd1608, -32'd1867, 32'd5969},
{32'd2925, 32'd1460, 32'd3991, 32'd440},
{32'd469, -32'd13963, -32'd6040, 32'd1286},
{32'd9919, 32'd10548, 32'd2283, 32'd8956},
{32'd10857, -32'd551, -32'd859, 32'd3006},
{32'd1050, -32'd5612, -32'd2132, -32'd4471},
{32'd6728, -32'd2184, 32'd2074, 32'd1158},
{32'd2824, -32'd2212, -32'd980, -32'd2968},
{32'd4594, -32'd4898, -32'd3692, 32'd7107},
{32'd10971, 32'd9887, 32'd3274, -32'd2115},
{32'd9528, 32'd1640, -32'd7007, -32'd1899},
{-32'd2398, 32'd2867, 32'd505, 32'd3137},
{-32'd5877, -32'd9255, 32'd4717, 32'd2425},
{32'd10623, 32'd5330, -32'd664, 32'd3427},
{32'd3820, -32'd5389, -32'd3939, -32'd1623},
{-32'd809, 32'd4503, 32'd6885, 32'd7432},
{-32'd13731, 32'd481, 32'd3515, -32'd6391},
{-32'd972, 32'd8752, 32'd7013, 32'd1057},
{-32'd3187, 32'd5084, 32'd882, 32'd3291},
{-32'd3831, -32'd299, -32'd1879, 32'd3907},
{-32'd9778, -32'd8956, 32'd1009, 32'd1562},
{-32'd13540, -32'd2337, 32'd3110, -32'd1212},
{-32'd327, 32'd5543, 32'd939, -32'd1768},
{32'd5225, -32'd5140, 32'd4184, -32'd7352},
{32'd8219, -32'd320, 32'd9118, 32'd8676},
{32'd17691, 32'd9905, -32'd3668, 32'd3480},
{-32'd2725, -32'd1699, 32'd7023, -32'd458}
},
{{32'd4769, 32'd9971, 32'd6981, -32'd1458},
{-32'd5185, -32'd5133, -32'd8898, -32'd8281},
{32'd3615, -32'd5096, -32'd1801, 32'd3975},
{-32'd44, 32'd1831, 32'd5758, 32'd1651},
{32'd3376, -32'd3670, 32'd7553, 32'd4353},
{32'd1224, -32'd11564, 32'd5449, -32'd9677},
{32'd13893, -32'd4031, -32'd20, -32'd3076},
{-32'd9612, -32'd2272, -32'd2800, 32'd3508},
{32'd5974, 32'd4585, -32'd1829, 32'd101},
{32'd7811, 32'd10962, 32'd2591, 32'd4703},
{-32'd11516, -32'd12969, 32'd847, 32'd6575},
{-32'd10456, -32'd10791, -32'd7384, 32'd6868},
{-32'd16323, 32'd4102, 32'd5887, 32'd4109},
{-32'd2611, 32'd18163, 32'd7944, 32'd7020},
{-32'd11247, -32'd4985, -32'd2953, 32'd10830},
{32'd785, 32'd3752, 32'd7801, 32'd7973},
{-32'd2965, 32'd11671, 32'd7618, 32'd875},
{-32'd8757, 32'd5869, 32'd466, 32'd4570},
{-32'd1111, 32'd379, 32'd1884, 32'd8216},
{-32'd3098, 32'd4578, 32'd6895, -32'd475},
{-32'd1563, -32'd5638, 32'd3024, -32'd149},
{32'd2613, -32'd13870, -32'd5746, -32'd2642},
{-32'd12156, -32'd908, -32'd3951, -32'd2039},
{-32'd1368, -32'd5105, -32'd6055, -32'd7591},
{32'd16238, -32'd3016, 32'd1551, 32'd5267},
{32'd7571, 32'd8598, 32'd8536, -32'd146},
{-32'd6049, 32'd3409, 32'd1666, 32'd4192},
{32'd9873, 32'd8756, -32'd1599, 32'd2141},
{-32'd796, 32'd3229, 32'd1060, -32'd2694},
{32'd5034, -32'd5165, -32'd8799, 32'd11752},
{32'd9614, 32'd1193, 32'd262, 32'd5073},
{-32'd2633, 32'd3685, -32'd1776, -32'd1809},
{32'd6184, 32'd4435, 32'd7090, 32'd3181},
{-32'd598, -32'd1652, -32'd6974, 32'd5375},
{32'd5974, 32'd10393, 32'd4703, 32'd2455},
{-32'd1326, -32'd8145, -32'd5926, 32'd12603},
{32'd628, -32'd3531, 32'd9829, -32'd3268},
{-32'd650, 32'd8727, 32'd12640, 32'd1001},
{32'd11434, 32'd7946, 32'd2089, 32'd2973},
{32'd750, -32'd1886, -32'd6859, 32'd1829},
{32'd5701, -32'd171, -32'd2944, -32'd8082},
{-32'd7710, -32'd6154, -32'd3402, 32'd9445},
{32'd654, 32'd11194, -32'd11544, -32'd1650},
{-32'd12671, -32'd3427, -32'd5517, 32'd6858},
{-32'd4771, -32'd10388, -32'd3766, -32'd128},
{-32'd7686, -32'd2085, -32'd5853, 32'd3964},
{-32'd16424, 32'd509, 32'd4816, 32'd4066},
{-32'd3353, -32'd3383, -32'd460, 32'd3020},
{-32'd1701, -32'd1008, -32'd7588, 32'd2608},
{32'd1885, 32'd2944, 32'd12334, -32'd6161},
{-32'd1821, -32'd2705, -32'd6890, -32'd589},
{-32'd1115, 32'd815, 32'd2695, -32'd4779},
{-32'd8779, 32'd8664, 32'd4982, 32'd5813},
{-32'd14360, 32'd11855, -32'd704, -32'd4190},
{-32'd5102, 32'd1443, -32'd100, 32'd11805},
{-32'd9238, -32'd12834, 32'd1041, -32'd8634},
{-32'd2506, 32'd3686, 32'd1707, -32'd356},
{32'd3033, -32'd9418, 32'd1139, -32'd9231},
{-32'd4063, -32'd2192, -32'd2739, -32'd10008},
{-32'd4530, 32'd7780, 32'd7265, -32'd4329},
{-32'd8679, -32'd216, -32'd1371, 32'd9305},
{32'd6403, -32'd2338, 32'd810, 32'd3668},
{-32'd10878, -32'd1087, -32'd3789, -32'd7828},
{-32'd9868, 32'd4605, 32'd2823, -32'd7140},
{-32'd4982, 32'd515, -32'd2187, 32'd14453},
{32'd8062, 32'd3136, 32'd3903, 32'd4316},
{-32'd1743, 32'd8374, 32'd6757, -32'd516},
{-32'd12566, -32'd8875, 32'd8392, 32'd923},
{-32'd2, 32'd2180, -32'd4537, 32'd3946},
{-32'd1057, -32'd6017, 32'd14454, -32'd6018},
{32'd1974, 32'd1146, 32'd2361, -32'd5951},
{32'd9485, -32'd772, 32'd6417, -32'd2154},
{32'd768, -32'd6613, 32'd1799, -32'd8062},
{-32'd3007, -32'd5207, -32'd4294, -32'd3106},
{32'd10192, -32'd423, 32'd4426, -32'd5465},
{-32'd12643, 32'd12871, 32'd6563, -32'd4818},
{-32'd12495, 32'd11718, -32'd2422, 32'd3310},
{-32'd6172, 32'd2707, 32'd8769, 32'd636},
{32'd11924, 32'd10912, -32'd1871, 32'd2488},
{-32'd1, 32'd2382, -32'd664, -32'd7729},
{32'd5399, 32'd1429, -32'd1718, -32'd1715},
{32'd3814, 32'd5800, -32'd5554, 32'd9392},
{32'd10196, -32'd468, -32'd1404, -32'd10830},
{32'd1133, 32'd13584, -32'd3842, -32'd4677},
{-32'd5858, -32'd7611, -32'd7087, 32'd4216},
{32'd11453, -32'd9867, -32'd5386, 32'd947},
{32'd2693, 32'd1280, 32'd9845, -32'd133},
{-32'd6265, -32'd6963, 32'd6113, -32'd7244},
{-32'd4185, -32'd3004, -32'd4871, 32'd1157},
{-32'd1640, -32'd5771, -32'd7231, -32'd941},
{32'd2179, -32'd3164, -32'd4731, 32'd2768},
{32'd3162, -32'd3779, -32'd6449, 32'd3172},
{-32'd2837, 32'd6312, -32'd8150, 32'd14119},
{32'd3553, 32'd8690, 32'd4364, 32'd60},
{-32'd15632, 32'd4670, 32'd4156, -32'd1457},
{-32'd2749, -32'd9721, -32'd1106, -32'd1539},
{32'd7212, 32'd10669, 32'd9318, 32'd1701},
{-32'd5458, -32'd469, 32'd5909, 32'd2672},
{-32'd10222, -32'd7727, -32'd2015, -32'd7163},
{32'd14979, 32'd7222, -32'd1003, 32'd909},
{-32'd9322, -32'd3349, 32'd6748, 32'd3109},
{-32'd4342, -32'd74, -32'd2519, -32'd713},
{-32'd11153, 32'd7339, -32'd590, 32'd2332},
{32'd16130, -32'd1051, -32'd939, 32'd5950},
{32'd1, -32'd10441, -32'd4508, 32'd706},
{32'd4564, -32'd5261, -32'd1132, 32'd5271},
{-32'd17086, 32'd1928, -32'd4667, -32'd7366},
{32'd7015, 32'd6385, -32'd3879, 32'd3847},
{-32'd8266, 32'd7210, -32'd9331, 32'd4062},
{-32'd22927, 32'd4677, 32'd1103, -32'd4293},
{32'd7845, -32'd3976, -32'd4414, -32'd1353},
{-32'd544, 32'd4045, -32'd4827, -32'd5558},
{32'd3099, 32'd7916, -32'd2228, 32'd2978},
{-32'd1555, -32'd2628, -32'd4371, -32'd7383},
{-32'd16387, 32'd4806, 32'd98, -32'd4589},
{-32'd15099, -32'd2964, 32'd2480, -32'd4606},
{32'd2090, -32'd5067, -32'd8850, -32'd8159},
{-32'd7109, 32'd3137, 32'd5207, -32'd1557},
{-32'd1795, -32'd1873, 32'd3135, 32'd5477},
{32'd11560, 32'd8401, 32'd10494, 32'd2513},
{-32'd5426, 32'd342, -32'd4729, 32'd2309},
{32'd8051, 32'd8607, 32'd6062, 32'd5241},
{32'd1287, 32'd6708, 32'd4162, 32'd2761},
{32'd2357, 32'd3234, 32'd3461, -32'd1677},
{-32'd849, -32'd9108, -32'd4408, 32'd8339},
{32'd35, 32'd7765, -32'd2910, -32'd914},
{-32'd7921, -32'd3686, -32'd10204, -32'd308},
{32'd9608, -32'd2376, -32'd7976, -32'd3776},
{-32'd3981, 32'd964, 32'd1693, 32'd893},
{32'd7033, -32'd373, -32'd409, -32'd8312},
{32'd1788, -32'd1260, -32'd296, -32'd11189},
{-32'd2054, 32'd918, -32'd873, -32'd3486},
{-32'd6797, -32'd7167, -32'd653, 32'd1078},
{32'd9868, -32'd4049, 32'd1151, 32'd211},
{32'd12984, 32'd6824, 32'd8182, -32'd6244},
{32'd930, -32'd3060, -32'd6934, -32'd6648},
{-32'd675, 32'd2630, -32'd2457, -32'd2720},
{-32'd2488, -32'd8940, 32'd5451, -32'd6941},
{-32'd2805, 32'd9422, 32'd3790, 32'd5500},
{-32'd11100, -32'd3409, 32'd2370, -32'd4351},
{32'd933, -32'd2097, 32'd2433, -32'd5321},
{-32'd3552, -32'd10210, -32'd4273, -32'd7645},
{32'd6520, 32'd3788, 32'd3544, -32'd504},
{-32'd6435, -32'd2363, -32'd4024, 32'd9646},
{32'd3929, -32'd2513, -32'd1161, 32'd12545},
{-32'd69, -32'd2805, -32'd7598, 32'd475},
{-32'd14158, 32'd1338, -32'd423, -32'd1366},
{-32'd2495, -32'd2643, -32'd13043, 32'd262},
{32'd812, -32'd116, 32'd12035, -32'd1542},
{-32'd14188, -32'd6704, 32'd1025, -32'd11112},
{-32'd8497, -32'd9823, -32'd6987, 32'd81},
{32'd13101, 32'd6020, -32'd6613, 32'd7739},
{-32'd17232, 32'd3742, -32'd4303, 32'd2257},
{-32'd9512, 32'd2328, 32'd9477, -32'd2455},
{-32'd10635, -32'd9861, -32'd7644, -32'd5318},
{-32'd447, -32'd696, 32'd1683, 32'd10504},
{-32'd5342, -32'd4351, 32'd4867, 32'd3103},
{32'd553, 32'd3655, 32'd4781, 32'd2683},
{32'd1667, -32'd1140, 32'd1997, -32'd156},
{-32'd7847, 32'd6297, -32'd10455, -32'd3160},
{32'd2925, 32'd2011, 32'd1587, 32'd4047},
{-32'd3187, 32'd6391, 32'd4839, 32'd3037},
{-32'd564, 32'd482, -32'd1235, -32'd8596},
{32'd20954, 32'd8769, -32'd7827, 32'd3356},
{-32'd2693, 32'd1631, 32'd558, 32'd2767},
{32'd4914, -32'd11113, 32'd4792, -32'd3305},
{-32'd1873, 32'd502, -32'd9052, 32'd8070},
{-32'd6365, -32'd10063, -32'd3860, -32'd2567},
{-32'd1828, 32'd5058, 32'd2848, 32'd272},
{-32'd4344, -32'd11550, 32'd8794, -32'd2736},
{-32'd4543, -32'd6085, -32'd8922, 32'd3918},
{-32'd3446, -32'd14620, 32'd398, -32'd3146},
{32'd6414, 32'd7181, 32'd8970, 32'd324},
{-32'd4227, -32'd9504, 32'd3799, 32'd10758},
{32'd1006, -32'd3861, 32'd1965, 32'd8046},
{32'd1368, 32'd6645, -32'd1673, 32'd4788},
{32'd1652, -32'd4579, -32'd634, 32'd1515},
{32'd1958, -32'd484, -32'd4226, -32'd11984},
{-32'd9605, 32'd15026, 32'd83, -32'd1699},
{-32'd621, -32'd9101, -32'd6611, -32'd1155},
{-32'd7541, -32'd4588, -32'd4942, 32'd2958},
{-32'd6914, 32'd1794, 32'd707, 32'd1184},
{-32'd7242, -32'd7614, 32'd4261, 32'd3430},
{-32'd5732, -32'd11149, -32'd3842, -32'd545},
{-32'd14298, -32'd8101, -32'd6248, 32'd10108},
{32'd20364, -32'd3772, 32'd4489, 32'd1103},
{32'd3571, 32'd2309, -32'd2386, 32'd503},
{32'd3980, -32'd2000, -32'd1209, -32'd3466},
{32'd2557, 32'd3481, -32'd3553, -32'd4661},
{32'd4061, -32'd131, -32'd7964, -32'd5598},
{-32'd12777, -32'd702, -32'd9951, 32'd3152},
{-32'd7357, 32'd3669, -32'd4182, 32'd4183},
{-32'd7087, 32'd976, 32'd3233, 32'd2527},
{32'd2393, -32'd890, -32'd2069, -32'd3626},
{32'd6405, 32'd7718, 32'd8638, -32'd5960},
{-32'd2884, -32'd7306, -32'd9780, 32'd992},
{32'd5305, -32'd5212, 32'd4200, 32'd114},
{32'd6285, 32'd2228, -32'd3481, 32'd415},
{32'd8389, -32'd3479, -32'd9812, 32'd1391},
{32'd2655, -32'd8583, 32'd6436, 32'd2978},
{-32'd3562, -32'd13622, -32'd4074, -32'd894},
{32'd12099, 32'd1628, -32'd3660, -32'd5603},
{32'd2724, -32'd10931, -32'd3306, -32'd4106},
{32'd2632, 32'd5645, 32'd4675, 32'd1425},
{32'd771, 32'd5229, -32'd7731, 32'd1610},
{-32'd6594, 32'd776, 32'd3132, -32'd10724},
{32'd15559, 32'd1046, -32'd347, 32'd8685},
{32'd3075, -32'd8361, -32'd3271, 32'd3652},
{32'd10830, 32'd11646, -32'd2046, -32'd1024},
{32'd11741, 32'd10220, 32'd4780, 32'd4264},
{32'd90, -32'd8232, 32'd5927, 32'd5955},
{32'd3328, 32'd3875, 32'd2892, 32'd4641},
{-32'd3011, -32'd4907, 32'd5296, -32'd5419},
{32'd8063, 32'd2289, 32'd2754, 32'd9415},
{-32'd10157, 32'd4396, -32'd474, -32'd8943},
{32'd10354, -32'd4541, -32'd9643, -32'd3711},
{-32'd1330, 32'd9447, 32'd10100, -32'd8461},
{32'd5160, -32'd4815, -32'd3382, 32'd1459},
{32'd3511, 32'd7126, 32'd8244, -32'd3273},
{-32'd1831, 32'd2228, -32'd7345, 32'd2311},
{32'd8338, 32'd6515, 32'd208, 32'd645},
{32'd1149, 32'd5377, 32'd3604, -32'd1850},
{32'd5113, 32'd3118, -32'd6490, -32'd4483},
{32'd4300, -32'd5753, 32'd2929, 32'd9839},
{-32'd22128, 32'd5860, -32'd903, 32'd1052},
{-32'd2501, -32'd12509, -32'd8359, -32'd2291},
{32'd9351, 32'd7701, -32'd9180, 32'd5813},
{32'd2810, -32'd10699, -32'd1406, 32'd3637},
{-32'd8733, 32'd496, 32'd776, -32'd3800},
{-32'd2729, 32'd10473, 32'd7826, -32'd11621},
{-32'd5224, 32'd6069, -32'd2669, -32'd6612},
{32'd5092, 32'd5900, -32'd4940, 32'd7670},
{32'd14296, -32'd11668, 32'd14872, -32'd5296},
{32'd6812, 32'd7172, -32'd10489, 32'd4161},
{-32'd805, -32'd202, 32'd1052, 32'd1043},
{-32'd6511, 32'd7168, 32'd2037, -32'd2527},
{32'd3534, -32'd5304, 32'd3691, 32'd10002},
{32'd8815, 32'd4026, 32'd9193, -32'd928},
{32'd2643, 32'd2419, 32'd6327, -32'd1707},
{32'd3364, 32'd3491, -32'd5571, -32'd3008},
{-32'd10396, 32'd855, 32'd6193, -32'd6752},
{32'd11080, 32'd3809, 32'd1817, -32'd169},
{-32'd6743, -32'd4272, -32'd5546, 32'd809},
{-32'd2596, 32'd2841, -32'd7084, 32'd5348},
{32'd483, 32'd13615, 32'd8185, -32'd714},
{32'd1522, 32'd4364, 32'd4473, 32'd1550},
{32'd6391, 32'd1603, -32'd11237, -32'd4024},
{32'd3441, -32'd2888, 32'd1131, 32'd394},
{-32'd3926, -32'd7335, -32'd4038, 32'd3489},
{32'd387, -32'd2402, 32'd6801, 32'd4651},
{-32'd8467, 32'd1775, -32'd12297, 32'd13605},
{32'd11704, 32'd11966, -32'd1730, 32'd3156},
{32'd6787, 32'd1757, 32'd6386, -32'd2440},
{32'd3654, 32'd4088, 32'd10887, 32'd4457},
{-32'd2983, 32'd5796, 32'd35, -32'd906},
{32'd11659, 32'd10454, 32'd5208, -32'd4394},
{32'd4261, -32'd17041, -32'd5770, 32'd3472},
{32'd6748, 32'd10411, -32'd1667, -32'd1366},
{32'd5687, -32'd13189, -32'd8196, 32'd2215},
{-32'd4394, 32'd4423, 32'd8788, 32'd2283},
{-32'd2413, -32'd7924, 32'd7647, 32'd5050},
{-32'd6863, 32'd7521, 32'd22, -32'd6526},
{-32'd1500, -32'd8163, 32'd4644, 32'd5447},
{32'd2259, -32'd6297, -32'd15605, -32'd6811},
{-32'd3331, -32'd11830, 32'd2563, 32'd8429},
{32'd11311, 32'd4374, -32'd3197, -32'd10063},
{32'd595, -32'd1709, -32'd1798, -32'd3533},
{32'd378, 32'd1547, -32'd7641, 32'd2362},
{-32'd7740, -32'd6612, -32'd5199, 32'd6028},
{-32'd671, 32'd1140, -32'd2006, -32'd21},
{32'd6502, -32'd189, 32'd8618, -32'd6379},
{32'd8557, -32'd4370, -32'd136, -32'd6132},
{-32'd7491, 32'd2811, -32'd8756, 32'd2502},
{-32'd1343, -32'd11004, -32'd2877, -32'd974},
{32'd6380, -32'd5140, 32'd6980, 32'd7642},
{-32'd7575, -32'd376, -32'd7118, -32'd3083},
{32'd5002, 32'd11278, 32'd3643, 32'd5497},
{-32'd2950, 32'd7136, -32'd2843, -32'd6412},
{32'd1704, -32'd10699, 32'd1761, 32'd1347},
{-32'd13322, -32'd26, -32'd6275, 32'd559},
{-32'd1136, 32'd7243, 32'd199, -32'd25},
{-32'd877, 32'd10209, -32'd5154, 32'd2046},
{-32'd10303, -32'd677, 32'd10470, -32'd335},
{32'd7781, 32'd6845, 32'd2395, -32'd3350},
{-32'd9321, -32'd6181, 32'd7573, 32'd3437},
{32'd893, -32'd1520, -32'd5434, -32'd4680},
{32'd9203, 32'd5602, -32'd4113, -32'd7507},
{-32'd4167, 32'd7029, 32'd5229, 32'd5028},
{32'd5517, 32'd7717, -32'd1980, 32'd2140},
{-32'd6207, 32'd1357, -32'd5848, -32'd4060},
{-32'd1459, 32'd1115, -32'd9408, 32'd880},
{32'd11803, -32'd2413, 32'd4547, -32'd1783},
{32'd3799, 32'd8463, -32'd7538, 32'd2341},
{32'd5481, -32'd4950, -32'd1757, 32'd2938},
{32'd10146, 32'd2483, -32'd2514, 32'd404},
{-32'd645, -32'd2099, -32'd2590, 32'd528},
{-32'd4851, 32'd8068, -32'd7813, 32'd9757},
{32'd6836, 32'd282, -32'd3894, -32'd742},
{32'd5913, 32'd140, -32'd1231, 32'd6356},
{32'd2111, -32'd7438, 32'd669, 32'd4021}
},
{{32'd10559, 32'd5626, 32'd4796, 32'd7087},
{-32'd5871, -32'd6774, -32'd7825, -32'd6789},
{32'd605, 32'd4069, 32'd1098, 32'd2031},
{-32'd1874, -32'd3221, 32'd1464, 32'd1360},
{-32'd2465, 32'd6610, 32'd2117, 32'd1384},
{-32'd1756, -32'd5230, -32'd5929, -32'd2616},
{-32'd2579, 32'd790, 32'd3982, 32'd4749},
{-32'd4412, -32'd1165, 32'd1286, -32'd2752},
{-32'd13600, -32'd444, 32'd2926, -32'd2937},
{32'd6982, 32'd13203, 32'd5570, 32'd3061},
{-32'd6214, 32'd3853, 32'd999, 32'd5089},
{32'd619, -32'd61, -32'd4194, 32'd2310},
{-32'd3379, 32'd9188, 32'd3243, 32'd2531},
{-32'd1367, -32'd4984, 32'd186, 32'd2186},
{-32'd19269, -32'd4354, 32'd2032, -32'd232},
{-32'd2911, -32'd2693, 32'd911, 32'd1545},
{32'd897, -32'd1230, -32'd3862, -32'd1461},
{32'd3512, 32'd359, 32'd1857, 32'd346},
{32'd1817, -32'd2788, -32'd7051, -32'd2815},
{32'd4057, 32'd3359, 32'd4467, 32'd3879},
{-32'd4171, 32'd582, -32'd205, 32'd63},
{32'd786, -32'd2650, -32'd5181, -32'd1699},
{-32'd5277, -32'd8847, -32'd307, -32'd10179},
{-32'd4192, -32'd5526, -32'd3744, -32'd2468},
{-32'd1935, 32'd3183, 32'd7332, 32'd2538},
{32'd4781, 32'd1971, -32'd569, 32'd9892},
{32'd9196, -32'd732, 32'd4427, -32'd5951},
{-32'd1468, 32'd3865, -32'd3803, -32'd4145},
{32'd3896, -32'd1556, -32'd6667, 32'd1912},
{-32'd1339, 32'd2023, 32'd2350, 32'd1306},
{-32'd2794, -32'd675, -32'd2257, 32'd4138},
{32'd1670, -32'd9358, -32'd7228, 32'd2602},
{32'd3637, 32'd3632, -32'd774, 32'd3398},
{-32'd9909, 32'd2832, -32'd1495, -32'd1919},
{32'd1612, 32'd9075, 32'd3608, 32'd2147},
{32'd667, -32'd7010, 32'd7664, 32'd1321},
{32'd1444, -32'd4213, 32'd389, -32'd2179},
{32'd7674, -32'd2161, -32'd6753, -32'd778},
{-32'd7586, 32'd6994, 32'd44, -32'd2925},
{32'd8468, -32'd8083, -32'd2438, -32'd1581},
{-32'd5964, 32'd3718, 32'd5690, -32'd6045},
{32'd6576, 32'd3021, 32'd6041, 32'd5269},
{32'd811, 32'd2762, -32'd5039, 32'd4626},
{-32'd10688, -32'd1119, 32'd529, -32'd5293},
{32'd8223, -32'd1837, -32'd4499, -32'd8425},
{32'd972, -32'd2077, 32'd5806, 32'd4872},
{32'd4608, 32'd655, -32'd4869, 32'd81},
{-32'd2453, -32'd7599, -32'd2670, -32'd2870},
{32'd4415, 32'd4568, 32'd2193, -32'd1131},
{32'd2007, -32'd1099, -32'd7161, 32'd3355},
{-32'd1685, -32'd6438, -32'd2003, -32'd5236},
{32'd1415, 32'd3716, 32'd3480, 32'd379},
{32'd14567, 32'd1556, -32'd4482, 32'd801},
{-32'd9932, 32'd161, -32'd3322, 32'd2223},
{-32'd9173, 32'd4470, -32'd2786, -32'd4971},
{-32'd3362, -32'd8352, 32'd765, -32'd4039},
{32'd6293, 32'd5316, 32'd815, -32'd6528},
{32'd2522, -32'd3324, -32'd114, -32'd646},
{-32'd4047, -32'd5684, -32'd6325, -32'd838},
{32'd8882, -32'd4324, -32'd5759, -32'd1604},
{-32'd8424, -32'd726, 32'd2735, -32'd2940},
{-32'd4210, 32'd2894, -32'd231, 32'd631},
{-32'd8324, -32'd9706, -32'd1584, -32'd3569},
{-32'd104, 32'd4291, 32'd2801, 32'd7654},
{32'd7426, -32'd1597, 32'd1100, -32'd4274},
{32'd8160, 32'd8833, -32'd696, 32'd7428},
{32'd663, -32'd5888, -32'd1351, -32'd2181},
{32'd14695, 32'd102, -32'd3198, -32'd6213},
{32'd2894, 32'd7053, 32'd5552, 32'd967},
{-32'd5257, -32'd5700, -32'd398, 32'd3912},
{32'd5256, 32'd5149, -32'd1115, 32'd965},
{32'd1716, 32'd2032, 32'd230, 32'd607},
{32'd14929, 32'd1629, -32'd1342, 32'd3881},
{-32'd3454, 32'd9138, 32'd3644, -32'd6107},
{-32'd1742, -32'd481, 32'd1701, 32'd6696},
{-32'd4123, 32'd4917, 32'd551, -32'd493},
{32'd2424, -32'd5334, -32'd190, -32'd1840},
{32'd3546, -32'd1821, -32'd2023, -32'd3996},
{-32'd1020, 32'd11274, 32'd7031, 32'd3742},
{32'd2059, -32'd1426, -32'd3430, -32'd3086},
{32'd1530, 32'd3087, 32'd3694, 32'd7511},
{32'd499, 32'd2420, -32'd610, -32'd1089},
{-32'd10256, -32'd2401, -32'd391, -32'd2852},
{-32'd5080, 32'd4479, -32'd7955, 32'd5010},
{-32'd489, 32'd4605, 32'd3689, -32'd7111},
{32'd132, -32'd8682, -32'd1905, -32'd229},
{-32'd805, 32'd6012, -32'd1370, 32'd1854},
{-32'd1594, -32'd4350, -32'd3381, -32'd6214},
{-32'd2906, 32'd3405, 32'd1927, -32'd6674},
{-32'd6607, 32'd1472, -32'd3731, -32'd3277},
{32'd8378, 32'd3376, 32'd8354, -32'd113},
{-32'd12330, -32'd5131, 32'd2867, -32'd1477},
{32'd8373, 32'd7068, -32'd562, 32'd8044},
{32'd4078, -32'd1770, 32'd3238, 32'd5832},
{32'd2246, -32'd2163, -32'd809, -32'd16},
{32'd5454, -32'd730, 32'd4192, 32'd1714},
{32'd7599, 32'd4198, 32'd6002, -32'd1599},
{-32'd1368, -32'd5979, 32'd3643, 32'd563},
{32'd663, 32'd3470, 32'd2665, 32'd3635},
{32'd8873, 32'd7453, 32'd2163, 32'd6495},
{32'd1877, -32'd5422, -32'd2936, 32'd2155},
{-32'd9208, 32'd2361, -32'd2163, 32'd547},
{32'd10721, -32'd1304, 32'd4814, -32'd4670},
{-32'd6515, 32'd8383, -32'd1389, -32'd1436},
{32'd3972, 32'd2332, 32'd3624, -32'd114},
{32'd5934, -32'd754, 32'd1248, 32'd7109},
{-32'd2871, -32'd12837, -32'd7351, 32'd5327},
{-32'd13190, -32'd4065, -32'd87, -32'd1064},
{-32'd2819, 32'd6519, 32'd4973, 32'd1919},
{32'd4599, -32'd1271, 32'd1948, 32'd1569},
{32'd142, 32'd9503, -32'd3054, -32'd5348},
{32'd8430, -32'd2668, 32'd3800, 32'd282},
{-32'd4097, -32'd27, 32'd1674, 32'd2623},
{32'd6476, -32'd4132, 32'd7428, 32'd1878},
{-32'd12937, 32'd450, 32'd1313, -32'd837},
{-32'd6889, -32'd1462, -32'd2544, -32'd5776},
{-32'd5099, 32'd2257, -32'd76, -32'd1989},
{-32'd3725, -32'd2411, 32'd3673, 32'd837},
{-32'd7245, -32'd2018, -32'd1088, -32'd1009},
{32'd526, 32'd10548, 32'd737, 32'd5020},
{-32'd2267, 32'd66, -32'd1451, -32'd3119},
{-32'd2736, 32'd5834, -32'd6572, -32'd2962},
{-32'd2865, 32'd5607, 32'd209, -32'd756},
{32'd6515, -32'd4594, -32'd1147, 32'd975},
{-32'd1630, -32'd2678, 32'd2912, -32'd365},
{-32'd1886, -32'd1861, -32'd3498, -32'd1119},
{-32'd918, -32'd7282, 32'd5015, -32'd6653},
{32'd1539, 32'd1845, -32'd1918, 32'd1289},
{32'd183, -32'd5878, -32'd2718, 32'd666},
{-32'd12139, 32'd2980, -32'd6821, -32'd5580},
{32'd7494, -32'd67, -32'd258, -32'd3017},
{32'd6353, -32'd2349, -32'd573, -32'd4409},
{-32'd1385, -32'd1888, -32'd1545, 32'd1136},
{32'd6628, 32'd2655, -32'd1310, -32'd1593},
{32'd2611, 32'd354, -32'd2090, 32'd1216},
{-32'd13161, 32'd1471, 32'd5577, 32'd644},
{-32'd6241, -32'd299, -32'd882, 32'd4675},
{32'd9046, -32'd1036, -32'd3142, 32'd4463},
{-32'd204, -32'd4618, 32'd6329, 32'd1330},
{-32'd3332, -32'd7032, -32'd2131, -32'd6226},
{32'd3355, -32'd2553, -32'd247, 32'd285},
{-32'd6386, -32'd2250, -32'd3701, -32'd352},
{-32'd1200, 32'd5669, -32'd2474, 32'd4752},
{-32'd1109, -32'd195, 32'd535, 32'd3787},
{-32'd3671, 32'd4688, 32'd1502, -32'd1067},
{-32'd5176, 32'd809, 32'd5459, 32'd3488},
{32'd754, 32'd300, -32'd1120, 32'd2},
{-32'd5756, -32'd8079, 32'd3016, 32'd3898},
{-32'd2396, 32'd1585, -32'd763, -32'd7115},
{32'd7056, -32'd5807, -32'd1712, -32'd5251},
{-32'd8321, -32'd2995, -32'd1566, -32'd1618},
{-32'd1712, -32'd2467, 32'd1260, 32'd4817},
{32'd2055, 32'd896, -32'd219, 32'd3154},
{-32'd4506, -32'd4429, -32'd2836, -32'd4161},
{-32'd8897, -32'd6858, -32'd1072, -32'd4339},
{-32'd2419, 32'd3836, -32'd2542, 32'd1072},
{32'd2193, 32'd5786, 32'd1410, 32'd10561},
{-32'd7702, -32'd1456, -32'd2047, 32'd1083},
{-32'd4395, -32'd2204, -32'd2701, -32'd1867},
{32'd10214, 32'd2985, 32'd7333, 32'd4425},
{32'd950, 32'd126, -32'd8671, 32'd293},
{32'd5224, 32'd4576, -32'd4024, -32'd3479},
{-32'd3931, -32'd3380, -32'd144, -32'd365},
{-32'd3471, 32'd8822, -32'd2941, 32'd4635},
{32'd5553, -32'd3179, 32'd1540, 32'd4606},
{-32'd3420, -32'd9967, -32'd908, -32'd2617},
{32'd3875, 32'd2609, -32'd8160, 32'd1907},
{-32'd6875, -32'd7208, -32'd2961, -32'd4477},
{-32'd5541, -32'd6295, -32'd3150, 32'd2504},
{32'd1712, -32'd5171, -32'd4074, -32'd4213},
{-32'd13098, -32'd4586, 32'd1100, -32'd1819},
{-32'd3177, -32'd4298, -32'd5112, -32'd925},
{32'd4732, 32'd9836, 32'd3729, 32'd7337},
{32'd671, -32'd872, -32'd2420, -32'd3868},
{-32'd3723, 32'd776, 32'd5818, 32'd7180},
{-32'd14334, 32'd8814, -32'd4040, -32'd7011},
{-32'd3959, -32'd3024, 32'd1467, -32'd3166},
{-32'd1585, 32'd919, -32'd1674, -32'd428},
{32'd1325, -32'd1813, 32'd4327, -32'd3110},
{-32'd9975, -32'd3303, -32'd5595, -32'd7263},
{-32'd7135, -32'd4567, 32'd3649, -32'd1927},
{32'd3094, -32'd3963, 32'd2662, -32'd5144},
{32'd4064, 32'd1285, 32'd311, -32'd2894},
{-32'd1261, 32'd2516, -32'd3553, -32'd2881},
{32'd851, 32'd3589, 32'd520, -32'd3502},
{-32'd807, 32'd7419, -32'd1209, -32'd832},
{32'd8161, -32'd275, 32'd539, 32'd8426},
{32'd426, 32'd5450, 32'd1573, -32'd1656},
{-32'd1929, 32'd6724, -32'd3485, 32'd4969},
{-32'd1426, -32'd4666, -32'd1983, 32'd501},
{-32'd7448, 32'd575, 32'd8169, 32'd852},
{32'd1118, -32'd6931, 32'd3060, 32'd1677},
{-32'd9543, -32'd1816, 32'd48, -32'd2358},
{32'd11630, -32'd10, -32'd4418, 32'd339},
{-32'd875, 32'd7509, 32'd3713, -32'd4047},
{32'd4560, -32'd866, 32'd3764, -32'd516},
{32'd4549, -32'd6639, -32'd219, 32'd6217},
{32'd78, -32'd2133, 32'd3392, 32'd356},
{-32'd11514, -32'd1053, -32'd8152, 32'd3929},
{32'd6346, 32'd4011, 32'd2238, -32'd2833},
{-32'd4904, -32'd9568, -32'd1322, -32'd1606},
{-32'd2883, 32'd1746, 32'd768, 32'd4219},
{32'd4661, 32'd2864, 32'd7959, -32'd1183},
{32'd10435, 32'd9, -32'd2453, 32'd3722},
{-32'd3221, -32'd6479, -32'd3806, -32'd7221},
{32'd17723, 32'd1703, 32'd215, 32'd1704},
{-32'd5981, 32'd8564, -32'd3288, 32'd1147},
{-32'd4810, 32'd1873, -32'd1001, -32'd7925},
{32'd959, 32'd950, 32'd1804, -32'd7767},
{32'd2437, 32'd4750, 32'd3166, 32'd236},
{32'd3428, -32'd4620, -32'd1334, -32'd5091},
{-32'd5686, 32'd5004, 32'd5081, -32'd3626},
{32'd787, -32'd4536, -32'd7491, 32'd3896},
{-32'd5943, 32'd3560, -32'd5567, 32'd794},
{32'd3037, 32'd5049, 32'd1894, -32'd517},
{-32'd7620, -32'd1118, -32'd2042, -32'd1857},
{-32'd2914, -32'd3083, -32'd3765, 32'd3703},
{-32'd14331, -32'd712, 32'd1397, 32'd3332},
{32'd8660, -32'd2582, 32'd2771, 32'd3254},
{32'd2398, 32'd4538, -32'd2240, 32'd3484},
{-32'd7839, 32'd164, -32'd3375, -32'd2889},
{-32'd1901, 32'd3978, 32'd5247, 32'd4381},
{32'd1673, 32'd3048, -32'd1903, -32'd85},
{32'd12307, -32'd2248, 32'd4132, -32'd1689},
{-32'd1695, 32'd2961, 32'd2138, 32'd5048},
{-32'd1413, 32'd5148, -32'd6276, -32'd445},
{-32'd892, -32'd5650, -32'd202, 32'd2288},
{32'd5965, -32'd1878, -32'd640, 32'd872},
{-32'd2670, 32'd558, 32'd397, 32'd246},
{32'd1512, -32'd3082, -32'd2078, -32'd4578},
{-32'd5255, 32'd3562, -32'd3421, 32'd143},
{-32'd279, -32'd2552, 32'd3070, -32'd2002},
{-32'd5455, -32'd3839, 32'd4191, 32'd9804},
{32'd5870, 32'd3901, -32'd165, 32'd1922},
{-32'd3876, -32'd5006, -32'd1907, -32'd4446},
{32'd1300, 32'd2883, 32'd3546, -32'd4616},
{-32'd6066, -32'd1605, -32'd2966, -32'd10153},
{-32'd2273, 32'd3510, -32'd3053, 32'd1727},
{32'd2629, -32'd1152, -32'd272, 32'd3057},
{-32'd20087, -32'd4044, 32'd443, -32'd5346},
{32'd2349, 32'd3984, 32'd1328, 32'd2497},
{-32'd4301, 32'd2686, 32'd1099, 32'd1524},
{-32'd13578, -32'd5821, 32'd796, -32'd2348},
{-32'd6604, -32'd4590, -32'd3054, 32'd2397},
{32'd1402, 32'd11953, 32'd8961, 32'd2048},
{32'd8998, 32'd599, -32'd6408, -32'd3014},
{-32'd5654, -32'd5854, -32'd3400, -32'd2849},
{-32'd762, -32'd2471, -32'd83, -32'd1238},
{-32'd3408, -32'd1313, -32'd3174, 32'd515},
{-32'd10536, -32'd963, 32'd1873, -32'd691},
{-32'd8384, 32'd3980, 32'd1432, 32'd2816},
{-32'd5216, 32'd1851, -32'd908, -32'd3278},
{32'd3541, 32'd8152, 32'd3175, -32'd6800},
{-32'd1495, -32'd713, -32'd884, 32'd9284},
{-32'd6077, 32'd270, 32'd487, 32'd1242},
{32'd1171, -32'd5891, -32'd1432, 32'd4088},
{-32'd5668, 32'd1770, -32'd438, -32'd6458},
{32'd4881, 32'd4211, 32'd8201, -32'd7228},
{-32'd6791, -32'd2550, -32'd3058, -32'd8334},
{32'd10156, 32'd4458, 32'd1133, -32'd2626},
{32'd3177, -32'd6348, -32'd3680, 32'd1859},
{-32'd186, 32'd6905, -32'd8855, 32'd1134},
{-32'd5140, -32'd4808, -32'd2182, -32'd965},
{32'd1661, 32'd4027, 32'd2231, -32'd1520},
{32'd5958, 32'd8098, -32'd1415, -32'd4832},
{32'd903, -32'd5400, 32'd706, -32'd935},
{32'd6822, 32'd3398, 32'd2135, 32'd2272},
{32'd2061, -32'd10365, 32'd1590, -32'd962},
{-32'd8866, -32'd5563, -32'd6474, -32'd8635},
{-32'd11694, -32'd5437, 32'd1376, -32'd830},
{32'd3211, -32'd806, -32'd5357, 32'd3712},
{-32'd1062, -32'd1151, -32'd5665, -32'd302},
{-32'd438, 32'd148, 32'd3824, -32'd1832},
{-32'd3108, 32'd2188, -32'd10127, -32'd23},
{-32'd12111, 32'd3344, -32'd3267, -32'd4832},
{-32'd8545, -32'd10091, 32'd2340, 32'd3633},
{32'd7972, 32'd13803, 32'd4815, 32'd4802},
{32'd5145, -32'd418, 32'd2538, -32'd4614},
{-32'd2114, -32'd9025, -32'd3732, -32'd5753},
{-32'd3579, -32'd198, -32'd3076, -32'd3674},
{-32'd3781, 32'd8039, 32'd510, 32'd6121},
{32'd2754, 32'd6111, -32'd431, 32'd7144},
{32'd8757, -32'd1604, 32'd3664, 32'd8207},
{32'd67, -32'd7676, 32'd3439, 32'd8337},
{-32'd2671, 32'd1143, 32'd1421, -32'd885},
{-32'd3732, -32'd4336, -32'd934, -32'd2474},
{32'd5743, 32'd4809, -32'd1357, -32'd2914},
{-32'd3431, 32'd2788, -32'd2900, -32'd158},
{-32'd4269, 32'd3341, 32'd3142, 32'd1781},
{-32'd3169, 32'd121, -32'd278, 32'd180},
{-32'd1434, 32'd2000, 32'd6883, -32'd2754},
{32'd12093, 32'd6620, 32'd3516, 32'd216},
{-32'd2316, -32'd5048, -32'd6270, 32'd4110},
{32'd4420, 32'd176, 32'd5397, -32'd319},
{-32'd8146, -32'd1498, -32'd4874, -32'd3265},
{-32'd5761, -32'd2083, 32'd851, -32'd1421},
{-32'd14402, -32'd1175, 32'd3357, 32'd3036},
{32'd3012, 32'd5866, 32'd5366, 32'd6092},
{32'd7270, 32'd8338, 32'd1399, 32'd3512},
{-32'd5659, -32'd5068, 32'd1209, -32'd6810}
},
{{32'd3848, 32'd5263, 32'd3934, 32'd2221},
{-32'd6518, -32'd1507, 32'd8153, -32'd854},
{-32'd2983, -32'd1188, -32'd1590, 32'd10613},
{32'd3782, 32'd827, 32'd14045, 32'd157},
{32'd10986, -32'd4108, -32'd2820, 32'd2846},
{-32'd8464, 32'd335, -32'd1742, -32'd3190},
{-32'd5467, -32'd5868, -32'd487, 32'd582},
{-32'd983, -32'd11607, 32'd3576, -32'd381},
{32'd7396, -32'd1686, -32'd8273, -32'd1692},
{32'd6280, 32'd7835, 32'd10006, 32'd7615},
{-32'd6381, -32'd4122, 32'd1534, 32'd2727},
{-32'd4005, 32'd6575, -32'd10674, -32'd6626},
{-32'd6274, 32'd3518, -32'd14419, -32'd9364},
{-32'd3023, -32'd12357, 32'd4296, 32'd4269},
{-32'd338, -32'd11357, -32'd4705, -32'd5918},
{-32'd1859, -32'd3274, 32'd4117, -32'd7713},
{32'd10637, 32'd1133, 32'd10251, 32'd5379},
{32'd4921, -32'd1706, 32'd5058, 32'd6291},
{-32'd1330, 32'd3726, -32'd7299, -32'd4303},
{-32'd12833, 32'd6092, 32'd5644, -32'd7139},
{-32'd5975, 32'd1567, -32'd1664, -32'd279},
{-32'd9955, -32'd9650, -32'd641, -32'd7578},
{-32'd10486, -32'd4509, 32'd3976, -32'd6118},
{-32'd873, -32'd11735, -32'd385, -32'd2038},
{-32'd95, 32'd6976, 32'd1886, 32'd1145},
{-32'd10387, -32'd5127, 32'd2757, 32'd3328},
{-32'd481, 32'd4074, -32'd6186, -32'd5876},
{-32'd4080, 32'd3705, -32'd3602, 32'd7918},
{-32'd4701, 32'd3688, 32'd1519, 32'd3309},
{-32'd8224, -32'd14187, -32'd6215, -32'd3521},
{32'd1480, -32'd7955, -32'd8803, -32'd4707},
{32'd1516, -32'd11428, -32'd969, -32'd7381},
{32'd8773, 32'd8742, 32'd373, 32'd8597},
{32'd3887, -32'd6382, -32'd5056, -32'd556},
{32'd5751, 32'd1941, 32'd9369, 32'd5869},
{-32'd2049, 32'd2731, -32'd1815, -32'd1709},
{32'd3060, -32'd4607, 32'd3251, 32'd2832},
{32'd269, -32'd2432, 32'd5591, 32'd5087},
{-32'd1781, 32'd3738, 32'd3273, -32'd6468},
{32'd1933, 32'd738, 32'd8767, -32'd2992},
{32'd4068, 32'd5558, 32'd1594, -32'd6480},
{32'd8195, 32'd2176, 32'd5920, -32'd539},
{32'd8958, -32'd1333, 32'd7985, 32'd4708},
{-32'd1444, -32'd12045, -32'd188, -32'd2293},
{-32'd5122, -32'd470, -32'd4372, -32'd124},
{32'd3888, 32'd8853, -32'd1364, -32'd2476},
{-32'd5074, -32'd9417, 32'd3255, -32'd7123},
{-32'd6159, -32'd2377, -32'd3528, -32'd4325},
{-32'd9047, 32'd422, 32'd13023, 32'd4949},
{-32'd1656, -32'd4122, 32'd4876, 32'd10018},
{-32'd4416, -32'd1992, -32'd2808, -32'd3646},
{-32'd27, 32'd4074, 32'd9309, 32'd3384},
{32'd6952, -32'd1831, -32'd4674, 32'd2903},
{32'd1550, -32'd3573, 32'd89, 32'd3026},
{32'd2878, -32'd4830, 32'd305, -32'd6150},
{32'd114, 32'd2232, -32'd367, -32'd1701},
{32'd16154, 32'd5274, 32'd15824, 32'd3377},
{-32'd6064, -32'd12518, -32'd2274, 32'd6604},
{32'd4182, -32'd1613, -32'd5289, -32'd5945},
{32'd3405, 32'd6240, 32'd1750, 32'd1620},
{32'd15774, -32'd2838, -32'd10362, -32'd155},
{32'd944, -32'd2483, -32'd9898, -32'd3090},
{-32'd7360, -32'd7011, -32'd11859, -32'd7645},
{32'd2464, -32'd2784, -32'd251, -32'd1840},
{32'd2289, 32'd6888, 32'd3969, 32'd3975},
{-32'd470, 32'd4447, 32'd8135, 32'd8597},
{32'd2393, 32'd4746, -32'd7146, -32'd1920},
{-32'd2990, 32'd3190, 32'd5707, 32'd3497},
{32'd1013, -32'd2819, -32'd9484, -32'd5702},
{32'd12984, -32'd10396, -32'd844, 32'd1360},
{-32'd1089, -32'd24, -32'd12543, 32'd2094},
{-32'd6878, -32'd1235, 32'd7068, 32'd7419},
{-32'd5384, -32'd10135, -32'd6284, 32'd907},
{-32'd1611, 32'd3979, 32'd5586, 32'd656},
{-32'd1892, -32'd1471, 32'd3313, 32'd8774},
{32'd398, -32'd4860, 32'd3925, -32'd2276},
{-32'd7511, -32'd10732, -32'd2261, 32'd6000},
{-32'd10509, 32'd5925, -32'd1692, -32'd2815},
{32'd11891, 32'd5360, 32'd4954, 32'd9314},
{32'd1065, -32'd6441, 32'd12759, 32'd4106},
{32'd11477, 32'd11686, -32'd1557, 32'd7626},
{32'd10604, 32'd5794, -32'd2071, -32'd2286},
{32'd6895, 32'd11136, -32'd1740, -32'd1629},
{32'd15635, 32'd3061, -32'd4748, 32'd5083},
{-32'd1671, -32'd6826, -32'd7388, 32'd1490},
{32'd6589, -32'd1603, -32'd9605, -32'd9650},
{32'd13888, -32'd8996, 32'd2974, 32'd7022},
{-32'd2827, -32'd14663, 32'd526, -32'd6598},
{32'd7285, -32'd3616, -32'd323, -32'd5826},
{32'd5637, -32'd2824, -32'd5272, -32'd4382},
{-32'd6448, 32'd629, 32'd4743, 32'd2186},
{32'd5151, -32'd3267, -32'd5034, -32'd2994},
{-32'd17952, -32'd4707, 32'd9604, 32'd2555},
{32'd6508, 32'd1649, 32'd17777, 32'd7603},
{-32'd7279, 32'd12819, 32'd1052, -32'd1052},
{-32'd484, -32'd7131, -32'd1408, 32'd386},
{32'd2801, -32'd151, 32'd4074, 32'd5804},
{-32'd173, -32'd2961, -32'd736, 32'd4447},
{32'd3249, -32'd1530, -32'd483, 32'd1292},
{32'd6013, 32'd9837, 32'd14696, 32'd6183},
{-32'd4282, -32'd6755, 32'd2265, 32'd6405},
{32'd3963, -32'd8340, -32'd8811, -32'd7846},
{32'd8562, -32'd1888, 32'd1347, -32'd2025},
{32'd3777, 32'd5307, -32'd7750, 32'd5136},
{-32'd1047, -32'd652, 32'd1967, -32'd723},
{32'd74, -32'd5603, 32'd2061, -32'd3182},
{-32'd11236, -32'd10663, -32'd7113, 32'd579},
{-32'd5567, -32'd8659, -32'd8399, 32'd6083},
{32'd4344, -32'd805, -32'd1429, -32'd7200},
{32'd4330, -32'd246, -32'd6552, 32'd2581},
{-32'd669, 32'd1973, 32'd1253, 32'd2783},
{32'd13128, -32'd1105, 32'd1629, -32'd1771},
{32'd6651, 32'd203, 32'd4839, 32'd4273},
{32'd6754, 32'd6235, 32'd7828, 32'd3070},
{32'd145, -32'd373, -32'd5428, -32'd2791},
{-32'd2719, 32'd24, 32'd877, -32'd4922},
{-32'd552, 32'd2213, 32'd8004, 32'd3883},
{-32'd6180, -32'd234, 32'd6321, -32'd641},
{32'd16611, -32'd4133, 32'd1955, -32'd3964},
{-32'd3178, 32'd13734, 32'd6837, 32'd2229},
{-32'd7815, 32'd7535, 32'd7846, -32'd8265},
{32'd5800, 32'd882, 32'd381, 32'd2200},
{-32'd11335, 32'd1858, 32'd4529, 32'd3854},
{-32'd6784, 32'd3700, 32'd4051, -32'd3219},
{32'd10634, -32'd890, -32'd13549, -32'd3509},
{-32'd2035, 32'd10502, 32'd5986, 32'd7198},
{-32'd5232, 32'd10378, 32'd2603, -32'd7911},
{-32'd2649, -32'd5852, 32'd2745, -32'd6314},
{32'd5031, 32'd3353, -32'd3128, -32'd9466},
{-32'd7188, 32'd1405, -32'd3874, 32'd11121},
{-32'd4125, -32'd1636, -32'd2068, -32'd4961},
{-32'd1619, -32'd1608, 32'd421, 32'd355},
{-32'd1745, 32'd7747, -32'd16317, -32'd7322},
{-32'd5220, 32'd14077, 32'd493, 32'd11151},
{32'd5221, 32'd2159, -32'd5352, -32'd10568},
{32'd6565, 32'd10711, -32'd4530, -32'd8186},
{-32'd1195, 32'd1078, -32'd1146, -32'd90},
{-32'd10931, 32'd13836, -32'd7197, -32'd3643},
{32'd2542, 32'd9127, -32'd2286, -32'd1426},
{-32'd9227, 32'd4173, -32'd65, -32'd4657},
{-32'd9724, -32'd6444, -32'd407, 32'd11747},
{32'd3476, -32'd3860, 32'd409, -32'd6275},
{32'd6324, 32'd4702, -32'd1323, 32'd663},
{32'd387, -32'd6916, -32'd495, -32'd4184},
{32'd13712, -32'd4668, 32'd576, 32'd9825},
{32'd1735, 32'd16203, 32'd7526, 32'd6988},
{32'd1868, -32'd7664, 32'd7089, 32'd1403},
{32'd4531, -32'd16041, -32'd11059, -32'd10355},
{-32'd5403, 32'd6315, -32'd2965, 32'd1241},
{-32'd4886, -32'd1373, -32'd4113, -32'd6842},
{-32'd286, -32'd3075, -32'd6134, -32'd2730},
{32'd7454, 32'd10337, 32'd2931, 32'd5984},
{-32'd4671, 32'd9942, 32'd1431, -32'd1500},
{32'd11092, -32'd2508, 32'd553, -32'd424},
{-32'd2755, -32'd10273, -32'd14802, -32'd8265},
{32'd12261, -32'd6278, -32'd3306, -32'd7877},
{-32'd1776, 32'd4702, 32'd5257, 32'd2462},
{32'd10309, 32'd4985, -32'd4544, -32'd3081},
{32'd2661, -32'd1679, -32'd3558, -32'd1741},
{32'd9146, -32'd1906, 32'd2378, -32'd7010},
{-32'd1249, -32'd1886, 32'd2758, -32'd1722},
{-32'd2164, -32'd2187, 32'd8923, -32'd322},
{-32'd4736, -32'd2878, -32'd7462, -32'd10185},
{32'd10693, -32'd1822, 32'd4665, 32'd1482},
{32'd953, 32'd3607, 32'd1587, 32'd8282},
{-32'd3911, 32'd1496, -32'd649, -32'd353},
{-32'd12398, -32'd912, 32'd5145, 32'd2684},
{32'd3036, -32'd4664, -32'd8998, -32'd9566},
{32'd3223, 32'd3632, 32'd8540, 32'd1702},
{32'd2632, -32'd8676, -32'd13107, -32'd587},
{-32'd650, -32'd6416, -32'd23, 32'd7244},
{-32'd1673, -32'd4463, -32'd3388, 32'd4844},
{32'd3962, 32'd3117, 32'd10635, 32'd5298},
{-32'd4080, 32'd1348, -32'd3949, 32'd2907},
{32'd635, 32'd866, -32'd9148, -32'd1158},
{32'd2764, -32'd2083, -32'd848, 32'd511},
{32'd6209, -32'd5302, -32'd2356, 32'd1316},
{32'd8803, -32'd687, -32'd84, -32'd860},
{-32'd4275, 32'd65, 32'd8107, -32'd988},
{-32'd3971, 32'd11054, -32'd289, -32'd3068},
{-32'd10579, -32'd7995, -32'd6778, -32'd5591},
{32'd677, -32'd8153, 32'd3760, -32'd1795},
{-32'd4708, 32'd1102, -32'd5919, -32'd3374},
{-32'd5581, 32'd63, -32'd5120, -32'd3885},
{-32'd7706, -32'd6078, -32'd3803, 32'd2348},
{32'd5234, 32'd13286, 32'd5930, -32'd916},
{-32'd178, 32'd7360, 32'd2630, 32'd3620},
{32'd130, -32'd3363, 32'd1324, 32'd164},
{32'd943, -32'd5473, 32'd6614, -32'd4479},
{32'd9676, 32'd3537, 32'd303, -32'd3947},
{32'd11829, 32'd789, 32'd3421, -32'd434},
{-32'd12777, -32'd9523, -32'd1036, 32'd1023},
{32'd8286, -32'd2328, 32'd3822, 32'd1272},
{32'd11967, -32'd650, 32'd1679, -32'd1275},
{-32'd8478, 32'd6728, 32'd3901, 32'd1930},
{-32'd380, -32'd4269, 32'd224, 32'd943},
{32'd907, 32'd191, -32'd7335, 32'd6965},
{-32'd3075, 32'd8444, 32'd1329, -32'd331},
{32'd1738, -32'd1348, 32'd7544, 32'd7931},
{32'd5774, -32'd2893, -32'd1207, -32'd3669},
{-32'd7190, -32'd11881, -32'd9088, -32'd3421},
{32'd7924, 32'd5230, -32'd4004, -32'd7049},
{32'd1324, 32'd13751, 32'd9156, -32'd494},
{-32'd5599, 32'd6240, 32'd9455, 32'd6751},
{-32'd4532, -32'd4158, -32'd1159, 32'd1475},
{-32'd6530, 32'd1508, 32'd7479, -32'd1899},
{32'd3376, 32'd6880, 32'd3445, 32'd2193},
{-32'd2781, -32'd16084, -32'd1817, -32'd1550},
{32'd7998, -32'd232, 32'd9174, 32'd5339},
{32'd7203, 32'd11673, 32'd7319, -32'd1665},
{-32'd382, -32'd11468, -32'd7425, 32'd3665},
{-32'd2495, -32'd588, 32'd1123, 32'd3348},
{32'd6324, 32'd122, -32'd514, -32'd11058},
{-32'd1158, -32'd7027, 32'd700, 32'd340},
{-32'd6538, 32'd4281, -32'd5122, -32'd3222},
{-32'd1220, -32'd13339, -32'd1928, 32'd4153},
{-32'd321, -32'd13826, 32'd9487, -32'd3199},
{-32'd5897, -32'd9938, -32'd6258, -32'd1787},
{32'd4111, 32'd12834, 32'd1267, 32'd4131},
{-32'd2465, 32'd920, -32'd3195, -32'd3966},
{-32'd12683, 32'd1138, 32'd6772, 32'd3312},
{-32'd7516, 32'd1612, 32'd3807, 32'd2586},
{32'd6391, 32'd5752, 32'd1993, -32'd5401},
{-32'd8861, 32'd5218, -32'd10871, -32'd5551},
{32'd1668, 32'd8820, -32'd10517, -32'd6328},
{32'd9106, -32'd10046, 32'd6069, 32'd3906},
{32'd1415, 32'd6523, 32'd8232, 32'd1017},
{32'd2208, -32'd3553, -32'd2091, -32'd4074},
{32'd2132, 32'd4707, 32'd3585, 32'd5974},
{-32'd1020, 32'd10542, 32'd7716, -32'd4474},
{-32'd3007, -32'd4997, -32'd5244, -32'd3548},
{32'd7704, 32'd10105, -32'd8219, -32'd4088},
{32'd6928, 32'd7707, 32'd2251, 32'd4892},
{-32'd4218, 32'd2121, -32'd1327, -32'd1665},
{-32'd3223, -32'd2908, 32'd833, 32'd1757},
{-32'd8059, -32'd5516, -32'd5291, -32'd3050},
{32'd2582, -32'd2274, -32'd4610, 32'd900},
{-32'd2394, 32'd11102, -32'd6299, 32'd6005},
{32'd15484, 32'd8637, -32'd1592, 32'd2798},
{32'd5273, 32'd3310, -32'd4668, -32'd885},
{32'd14210, 32'd8266, 32'd1926, -32'd607},
{32'd3536, -32'd2804, -32'd4080, -32'd4149},
{32'd270, -32'd7380, -32'd1636, -32'd7870},
{32'd11947, 32'd4995, 32'd10185, 32'd9937},
{32'd11383, 32'd11703, 32'd8369, 32'd6960},
{32'd11311, 32'd2205, 32'd81, -32'd935},
{-32'd9459, -32'd1748, -32'd420, -32'd1836},
{-32'd8266, 32'd13111, 32'd635, -32'd1312},
{-32'd15009, 32'd3742, 32'd5294, -32'd126},
{32'd173, -32'd7434, -32'd4405, -32'd1314},
{32'd13174, -32'd3696, 32'd11277, -32'd4126},
{32'd1833, -32'd765, -32'd10453, 32'd8861},
{-32'd5918, 32'd11416, 32'd2418, 32'd4455},
{32'd1134, -32'd8430, -32'd525, 32'd1307},
{-32'd4919, -32'd3540, -32'd49, -32'd7181},
{32'd7094, 32'd4717, 32'd8315, 32'd739},
{32'd6790, 32'd4712, -32'd1092, -32'd3765},
{32'd533, 32'd8202, -32'd4248, -32'd3055},
{-32'd1073, -32'd5092, 32'd75, -32'd651},
{-32'd1249, 32'd12700, -32'd577, 32'd4692},
{-32'd2288, -32'd1799, 32'd6918, 32'd873},
{32'd13501, -32'd2753, -32'd3431, -32'd1351},
{-32'd3643, -32'd5155, 32'd1329, 32'd5645},
{-32'd6754, -32'd0, -32'd11659, -32'd2854},
{-32'd6975, 32'd1880, 32'd3945, 32'd7257},
{-32'd2498, -32'd1629, -32'd6819, 32'd1165},
{32'd13451, 32'd8262, -32'd5532, 32'd3153},
{32'd12605, 32'd2940, -32'd6054, -32'd4141},
{32'd6739, -32'd4696, 32'd3292, -32'd4823},
{32'd6083, 32'd4028, 32'd272, 32'd3939},
{-32'd9924, -32'd4779, -32'd6070, 32'd4192},
{-32'd5151, -32'd2201, 32'd5784, 32'd4011},
{-32'd11492, -32'd8232, -32'd3410, -32'd8263},
{-32'd8393, -32'd11894, -32'd6371, -32'd2547},
{-32'd2792, -32'd297, -32'd7291, -32'd582},
{-32'd4569, -32'd927, -32'd1403, 32'd3372},
{32'd11964, 32'd13145, 32'd10929, 32'd8223},
{-32'd12159, 32'd3160, -32'd5247, -32'd1413},
{-32'd2938, -32'd6466, -32'd11748, -32'd10036},
{32'd6879, -32'd1662, -32'd4505, -32'd5919},
{32'd9906, 32'd4004, 32'd8353, 32'd6839},
{32'd9901, 32'd7956, -32'd2688, 32'd1727},
{32'd4, 32'd9110, -32'd73, -32'd4976},
{-32'd8822, 32'd2699, 32'd6716, 32'd8089},
{32'd3097, 32'd7060, -32'd6221, -32'd1487},
{-32'd4382, -32'd7674, 32'd143, -32'd4169},
{32'd10615, 32'd4947, 32'd1324, 32'd2646},
{-32'd4685, -32'd7490, 32'd7376, -32'd1322},
{32'd2070, -32'd6465, -32'd5233, 32'd6771},
{32'd3064, 32'd2704, 32'd5875, -32'd1107},
{-32'd474, -32'd3354, 32'd3922, -32'd5944},
{32'd7914, 32'd2121, 32'd5462, 32'd3790},
{32'd12074, 32'd10414, 32'd6007, 32'd3733},
{-32'd12816, 32'd1838, -32'd4628, -32'd5634},
{-32'd11476, -32'd8075, -32'd9825, -32'd5818},
{-32'd11128, -32'd14748, -32'd5061, -32'd713},
{32'd10779, -32'd4135, 32'd4480, 32'd4581},
{-32'd2388, -32'd7936, -32'd3150, -32'd2250},
{32'd8513, -32'd3865, 32'd9277, -32'd745},
{-32'd4728, 32'd2131, -32'd3905, -32'd5863}
},
{{32'd6239, -32'd4185, 32'd2944, -32'd1384},
{32'd5039, -32'd9631, -32'd4265, -32'd297},
{32'd9353, 32'd5418, -32'd1625, -32'd4888},
{-32'd3424, 32'd2254, 32'd4423, 32'd5651},
{-32'd4363, 32'd7084, 32'd1607, -32'd6101},
{32'd9246, -32'd3848, 32'd2209, 32'd708},
{-32'd1462, -32'd5341, -32'd23, 32'd2869},
{32'd1459, -32'd10165, -32'd8996, 32'd5375},
{-32'd1570, 32'd259, -32'd1754, 32'd767},
{32'd5203, 32'd7347, 32'd5821, 32'd7146},
{-32'd10294, 32'd1894, 32'd13475, 32'd3394},
{-32'd8275, 32'd34, -32'd2952, -32'd12059},
{-32'd2423, -32'd1113, -32'd1335, -32'd1335},
{32'd3361, -32'd7976, -32'd800, -32'd6916},
{-32'd4727, -32'd6436, 32'd1276, -32'd730},
{32'd3950, -32'd3480, -32'd6264, -32'd12421},
{32'd2909, 32'd6909, -32'd361, -32'd8752},
{32'd8244, -32'd3903, -32'd6495, -32'd5544},
{32'd5451, 32'd1503, -32'd2588, 32'd13126},
{-32'd8830, 32'd8476, 32'd4245, -32'd4586},
{32'd11144, 32'd11901, 32'd3773, 32'd1379},
{-32'd3433, -32'd2277, -32'd7992, 32'd9049},
{-32'd2450, -32'd1319, 32'd2604, 32'd7931},
{-32'd5264, -32'd2783, 32'd842, -32'd1211},
{32'd13013, 32'd3851, 32'd731, 32'd1720},
{32'd6357, 32'd9325, -32'd2939, 32'd4905},
{-32'd8464, 32'd667, 32'd2849, 32'd372},
{32'd3634, 32'd2355, -32'd289, 32'd1006},
{-32'd1222, -32'd552, 32'd413, -32'd1675},
{-32'd623, 32'd6329, 32'd237, -32'd1293},
{-32'd1254, -32'd3121, 32'd4229, 32'd1926},
{-32'd5289, -32'd1991, 32'd3222, -32'd8727},
{32'd6981, 32'd2304, 32'd367, -32'd3166},
{32'd262, -32'd3707, -32'd7424, 32'd2470},
{32'd3350, 32'd1699, 32'd5747, 32'd9089},
{-32'd4865, -32'd3005, 32'd4443, -32'd10222},
{32'd12636, 32'd4680, -32'd9516, -32'd978},
{32'd11072, -32'd6089, -32'd549, -32'd5599},
{-32'd3477, -32'd3711, -32'd72, 32'd1469},
{32'd4884, -32'd1273, 32'd2408, -32'd3149},
{-32'd1841, 32'd10522, 32'd8526, 32'd12975},
{-32'd3554, 32'd6604, 32'd6981, 32'd716},
{-32'd12015, 32'd1399, 32'd2890, 32'd3275},
{32'd6163, 32'd1213, -32'd16121, 32'd871},
{32'd1109, -32'd17537, -32'd5180, -32'd1847},
{32'd12848, -32'd13665, 32'd2552, -32'd3823},
{-32'd3383, -32'd4563, 32'd2268, 32'd2183},
{32'd1186, -32'd17120, -32'd10565, -32'd10333},
{32'd4844, -32'd559, 32'd567, -32'd1009},
{-32'd1513, -32'd1172, -32'd3124, -32'd511},
{-32'd15922, 32'd1752, -32'd1236, -32'd12045},
{-32'd6955, 32'd2353, -32'd630, 32'd3905},
{-32'd750, 32'd7392, -32'd3467, -32'd6866},
{-32'd13260, -32'd6432, 32'd3454, 32'd5662},
{32'd2250, -32'd588, -32'd59, 32'd987},
{32'd6130, -32'd9506, -32'd2609, -32'd5562},
{32'd895, -32'd743, -32'd13766, 32'd2114},
{32'd2749, -32'd160, -32'd2900, -32'd3802},
{32'd2629, -32'd3132, 32'd125, -32'd1430},
{-32'd2227, -32'd7536, 32'd5088, -32'd10334},
{32'd1311, 32'd7946, -32'd6950, -32'd9186},
{32'd13409, -32'd1853, 32'd1153, -32'd5495},
{-32'd10099, -32'd3092, 32'd17644, -32'd4004},
{32'd4722, -32'd8071, -32'd3149, -32'd3438},
{-32'd926, -32'd3151, 32'd2420, 32'd3452},
{32'd5100, 32'd9722, 32'd11570, -32'd2814},
{-32'd676, 32'd2006, -32'd2370, 32'd5178},
{-32'd200, -32'd763, 32'd10067, -32'd12097},
{-32'd11085, -32'd3559, -32'd9524, -32'd1529},
{32'd8450, -32'd12767, 32'd4078, 32'd3466},
{32'd9353, -32'd4412, 32'd5202, -32'd251},
{32'd16117, -32'd8725, -32'd2646, 32'd5925},
{32'd6919, -32'd387, -32'd5650, -32'd5573},
{-32'd9108, 32'd3448, -32'd3042, -32'd171},
{32'd3542, 32'd5597, -32'd3552, 32'd2518},
{32'd4957, -32'd2828, -32'd8988, 32'd2898},
{32'd1233, -32'd1358, -32'd5879, 32'd1355},
{-32'd1812, -32'd3029, -32'd4402, -32'd2010},
{32'd18670, 32'd5175, 32'd9858, 32'd98},
{-32'd12740, 32'd11912, -32'd10514, -32'd6442},
{32'd2021, 32'd3419, 32'd9920, 32'd4387},
{32'd697, 32'd5509, 32'd11074, 32'd6556},
{-32'd1832, -32'd8053, -32'd1263, 32'd3977},
{32'd6698, -32'd10611, 32'd13735, 32'd4755},
{-32'd9283, 32'd3018, -32'd9384, -32'd19349},
{-32'd681, 32'd1035, 32'd4727, 32'd2941},
{32'd5271, 32'd5099, 32'd5627, -32'd953},
{-32'd9510, -32'd9802, -32'd972, -32'd3396},
{-32'd1788, 32'd1449, -32'd8698, -32'd358},
{-32'd1873, -32'd10041, -32'd3461, -32'd546},
{-32'd2488, 32'd128, 32'd3435, -32'd1629},
{32'd4750, -32'd8205, 32'd4525, -32'd12317},
{32'd3328, 32'd7837, 32'd923, -32'd1992},
{-32'd863, 32'd3791, 32'd6458, 32'd6397},
{32'd1577, 32'd9869, 32'd1454, -32'd4165},
{32'd4111, -32'd7808, 32'd9048, 32'd537},
{-32'd2770, 32'd8450, 32'd5167, 32'd1713},
{32'd7260, -32'd5856, -32'd13199, -32'd1652},
{-32'd1928, 32'd6864, -32'd4182, -32'd9822},
{32'd6929, -32'd753, 32'd2335, -32'd2091},
{32'd3133, -32'd4889, -32'd97, -32'd562},
{32'd1248, -32'd4718, 32'd10394, 32'd2728},
{32'd2626, 32'd5965, 32'd5482, 32'd9051},
{32'd13298, 32'd4205, 32'd6523, 32'd2369},
{32'd1202, 32'd5813, -32'd6625, -32'd1137},
{32'd6277, 32'd6688, 32'd8920, 32'd2273},
{-32'd2628, -32'd4347, 32'd1886, 32'd7990},
{-32'd11645, -32'd307, -32'd76, 32'd361},
{-32'd1433, 32'd9069, 32'd10364, 32'd4178},
{-32'd4607, -32'd12896, -32'd3513, -32'd8435},
{-32'd5572, -32'd7337, -32'd2508, -32'd1931},
{-32'd1812, -32'd205, 32'd2288, -32'd2339},
{32'd1415, 32'd2881, -32'd2501, 32'd7443},
{-32'd858, 32'd12246, 32'd9535, -32'd4745},
{-32'd3248, 32'd1950, 32'd3161, 32'd7783},
{-32'd2215, 32'd339, 32'd2610, -32'd8336},
{-32'd8434, 32'd4893, -32'd3184, 32'd6221},
{32'd3155, 32'd1369, -32'd7929, 32'd3835},
{32'd10428, -32'd1821, 32'd10613, 32'd9371},
{32'd11245, 32'd7756, 32'd5822, -32'd766},
{-32'd4902, 32'd11379, -32'd1073, 32'd1779},
{32'd797, 32'd3979, -32'd2741, -32'd2965},
{-32'd6022, -32'd10379, -32'd15402, -32'd4223},
{32'd4148, 32'd9759, 32'd2800, 32'd2389},
{-32'd7683, -32'd167, -32'd7734, -32'd4539},
{32'd19660, 32'd3844, 32'd924, -32'd1362},
{32'd3411, 32'd258, 32'd175, -32'd1716},
{-32'd3902, 32'd7585, -32'd4129, 32'd2119},
{-32'd18195, -32'd4908, -32'd6403, 32'd3503},
{32'd5788, -32'd228, -32'd9120, -32'd8213},
{-32'd13573, -32'd9140, -32'd12317, -32'd1327},
{-32'd7080, -32'd7937, 32'd26, 32'd115},
{-32'd3140, -32'd11926, 32'd380, -32'd2027},
{-32'd223, 32'd6038, -32'd6822, 32'd4373},
{-32'd7871, 32'd5257, -32'd6009, -32'd584},
{-32'd10043, -32'd4216, 32'd3448, -32'd9562},
{32'd6913, 32'd3478, 32'd6075, -32'd104},
{-32'd10175, 32'd2811, 32'd6820, -32'd2041},
{-32'd4559, 32'd14853, 32'd448, -32'd7808},
{-32'd7541, -32'd18877, -32'd10009, -32'd4136},
{-32'd11249, -32'd7277, -32'd1237, 32'd5551},
{32'd1563, -32'd7883, 32'd5877, 32'd9780},
{32'd1819, 32'd12220, 32'd2491, -32'd8224},
{-32'd8676, -32'd6093, 32'd3798, -32'd1108},
{32'd17454, -32'd79, 32'd4197, -32'd4521},
{-32'd3881, 32'd7673, -32'd5479, 32'd1417},
{-32'd534, -32'd1209, -32'd4050, 32'd2959},
{32'd2891, -32'd6928, -32'd9902, 32'd344},
{32'd9013, 32'd1384, 32'd6789, -32'd1786},
{-32'd7905, -32'd4496, -32'd3074, -32'd576},
{-32'd6415, -32'd5273, -32'd3904, -32'd1328},
{-32'd1782, 32'd2445, 32'd13609, 32'd2633},
{-32'd1178, -32'd6919, -32'd1624, -32'd12824},
{-32'd3716, 32'd3190, -32'd1337, 32'd708},
{-32'd12562, -32'd14360, 32'd1899, -32'd6084},
{-32'd6104, 32'd77, -32'd9153, 32'd8268},
{32'd409, 32'd9329, 32'd5575, 32'd7390},
{-32'd4616, -32'd5173, -32'd10, 32'd430},
{32'd2092, 32'd1103, 32'd5341, 32'd5892},
{-32'd6395, 32'd3904, -32'd3455, -32'd8453},
{-32'd10849, -32'd2713, 32'd1363, 32'd2085},
{32'd5969, 32'd1774, -32'd5357, 32'd566},
{-32'd6633, 32'd2652, 32'd2764, 32'd1095},
{-32'd1569, 32'd8299, 32'd9243, 32'd7776},
{32'd17658, 32'd9102, -32'd1745, -32'd2702},
{32'd2848, -32'd7454, 32'd1224, 32'd5956},
{32'd5633, -32'd846, 32'd6335, 32'd10924},
{-32'd7934, 32'd462, -32'd7628, -32'd5492},
{-32'd2049, -32'd11623, -32'd3484, -32'd8571},
{-32'd6177, -32'd7863, -32'd3182, -32'd3848},
{32'd1791, -32'd9710, 32'd281, -32'd6503},
{-32'd4101, -32'd4179, -32'd1865, 32'd486},
{32'd2708, 32'd2954, 32'd15944, 32'd1832},
{32'd4219, -32'd2673, 32'd1947, 32'd6277},
{32'd13918, 32'd11189, 32'd8200, 32'd1217},
{32'd680, 32'd3308, -32'd370, 32'd4294},
{32'd8722, 32'd328, 32'd10279, 32'd4226},
{32'd10347, -32'd5334, -32'd1833, -32'd3934},
{-32'd3733, 32'd10564, 32'd7281, -32'd643},
{32'd674, -32'd5415, -32'd11901, 32'd4075},
{-32'd3249, 32'd250, 32'd3478, 32'd1155},
{-32'd5765, -32'd17714, -32'd579, -32'd96},
{32'd3386, 32'd3328, 32'd691, -32'd4422},
{-32'd7628, -32'd2247, 32'd9019, -32'd3299},
{32'd4585, 32'd6947, 32'd15097, 32'd9057},
{32'd17253, 32'd3907, 32'd2966, -32'd3091},
{-32'd1280, 32'd1471, 32'd7352, -32'd147},
{-32'd9725, 32'd2149, 32'd7483, -32'd6034},
{32'd2374, 32'd2321, 32'd6784, -32'd4900},
{-32'd13065, 32'd3402, 32'd5326, 32'd12013},
{32'd10238, 32'd4969, -32'd305, -32'd5030},
{32'd1441, -32'd5236, -32'd1971, -32'd1360},
{32'd14562, -32'd12112, 32'd2184, 32'd5425},
{32'd2723, 32'd10194, 32'd232, -32'd4344},
{32'd2237, -32'd14022, -32'd4766, -32'd15438},
{-32'd7155, 32'd321, -32'd5651, 32'd1642},
{32'd749, 32'd9882, 32'd5301, -32'd3696},
{32'd6315, 32'd337, -32'd1036, -32'd2824},
{-32'd4558, -32'd11375, 32'd651, 32'd2762},
{32'd4729, -32'd1113, -32'd2097, 32'd2212},
{-32'd8390, -32'd13055, -32'd4938, -32'd1335},
{-32'd7192, -32'd3187, 32'd6920, 32'd11439},
{-32'd2791, -32'd4775, -32'd6547, -32'd858},
{-32'd4148, 32'd1645, 32'd2870, 32'd3244},
{-32'd1509, -32'd2992, -32'd12230, -32'd323},
{-32'd8726, -32'd4901, -32'd266, 32'd5409},
{32'd2495, 32'd1052, -32'd61, -32'd2010},
{-32'd9368, 32'd3594, -32'd4717, -32'd10621},
{32'd7607, -32'd7626, -32'd1496, 32'd8409},
{-32'd10866, 32'd4200, -32'd9102, -32'd9930},
{32'd1751, -32'd5714, -32'd522, -32'd417},
{32'd7507, -32'd9528, 32'd4333, -32'd2361},
{-32'd2987, 32'd4893, 32'd17005, -32'd2113},
{32'd11832, -32'd6086, -32'd7046, -32'd1554},
{-32'd6541, -32'd1217, 32'd4198, 32'd6525},
{32'd771, -32'd7781, -32'd1350, 32'd7551},
{-32'd624, -32'd6416, 32'd5349, 32'd3433},
{-32'd1095, 32'd1350, 32'd4167, 32'd7664},
{32'd2769, 32'd857, 32'd1440, 32'd7391},
{32'd6627, 32'd13649, -32'd182, 32'd4851},
{-32'd4696, -32'd105, 32'd6046, -32'd1007},
{-32'd5007, 32'd12607, 32'd9447, 32'd1344},
{32'd17257, 32'd8646, -32'd663, -32'd1726},
{-32'd2449, 32'd5934, -32'd3612, 32'd81},
{-32'd7931, 32'd5356, -32'd3970, -32'd6057},
{32'd1870, -32'd601, -32'd6126, 32'd877},
{-32'd5868, 32'd3733, -32'd6084, 32'd15074},
{32'd8486, -32'd4136, -32'd7746, 32'd2609},
{-32'd17811, -32'd12085, -32'd8537, 32'd7067},
{-32'd3470, 32'd7476, 32'd676, 32'd890},
{-32'd12055, -32'd13502, 32'd7233, 32'd1266},
{-32'd8287, -32'd5164, -32'd2712, -32'd991},
{32'd6477, 32'd4251, 32'd4654, -32'd3558},
{-32'd14925, 32'd5943, -32'd1257, -32'd1327},
{32'd2899, -32'd1796, 32'd1010, 32'd10525},
{32'd4206, -32'd12763, -32'd3654, -32'd3861},
{-32'd795, -32'd7431, -32'd4632, -32'd3185},
{32'd8940, -32'd2534, 32'd11082, -32'd2131},
{32'd113, 32'd8847, 32'd14256, 32'd902},
{-32'd563, -32'd4789, -32'd13793, -32'd5892},
{-32'd5220, 32'd13622, -32'd499, -32'd4199},
{32'd560, 32'd8211, 32'd2003, -32'd9551},
{-32'd4326, -32'd2556, -32'd6756, 32'd5518},
{32'd12747, 32'd6252, 32'd6435, -32'd6246},
{32'd8969, 32'd3969, 32'd11750, 32'd3413},
{-32'd2915, 32'd6396, -32'd13637, -32'd214},
{-32'd12165, -32'd9005, 32'd2719, -32'd3488},
{32'd10088, -32'd228, 32'd4808, -32'd4491},
{32'd3722, 32'd3658, -32'd369, 32'd12074},
{32'd14893, -32'd1772, 32'd8580, 32'd4470},
{32'd376, 32'd5672, 32'd2303, -32'd5961},
{-32'd10498, -32'd6336, -32'd3828, 32'd4591},
{32'd7649, 32'd5173, -32'd6148, -32'd6150},
{-32'd3879, -32'd117, 32'd15755, 32'd12208},
{-32'd15187, 32'd5833, 32'd1983, 32'd5790},
{-32'd5219, -32'd12444, 32'd4649, 32'd13156},
{-32'd4485, 32'd5353, 32'd7300, 32'd4411},
{-32'd8990, 32'd2028, 32'd435, 32'd3988},
{-32'd24894, -32'd8501, 32'd5489, 32'd7060},
{32'd10432, -32'd4920, 32'd8661, -32'd8570},
{32'd4548, -32'd6948, 32'd4380, -32'd445},
{32'd8148, 32'd9624, 32'd6133, -32'd1402},
{32'd6273, -32'd12718, -32'd6197, -32'd3766},
{32'd7943, -32'd7958, -32'd6021, -32'd4309},
{32'd7738, -32'd1194, 32'd22, 32'd4493},
{32'd7249, 32'd4787, 32'd2305, -32'd13762},
{-32'd3327, 32'd12071, 32'd4483, 32'd1918},
{-32'd7009, 32'd4817, -32'd1028, -32'd9664},
{32'd2872, -32'd9244, -32'd627, 32'd3088},
{32'd1368, -32'd6518, -32'd2296, 32'd645},
{32'd9198, 32'd333, 32'd7727, 32'd648},
{32'd10308, 32'd3265, -32'd7771, 32'd1025},
{32'd8961, -32'd3349, 32'd813, 32'd2572},
{32'd9843, -32'd11292, -32'd2586, -32'd5617},
{32'd4946, 32'd10119, 32'd11602, 32'd2613},
{32'd1087, -32'd7957, -32'd7499, 32'd4463},
{32'd4297, 32'd5674, 32'd3465, 32'd1657},
{32'd7633, 32'd12563, 32'd640, -32'd7388},
{32'd7022, 32'd3613, -32'd14734, 32'd1207},
{-32'd5192, 32'd503, -32'd3737, -32'd6557},
{32'd9487, 32'd4362, -32'd2658, 32'd4508},
{32'd5656, 32'd2065, 32'd13683, -32'd6669},
{-32'd14799, -32'd5880, 32'd7849, -32'd690},
{32'd3116, -32'd1344, 32'd3144, 32'd3726},
{-32'd3435, -32'd753, 32'd7725, -32'd3308},
{-32'd11641, -32'd11196, -32'd3331, 32'd2073},
{32'd7580, 32'd3494, -32'd1499, 32'd2597},
{32'd4949, 32'd1601, -32'd7099, -32'd3410},
{-32'd3009, 32'd1985, -32'd2307, -32'd8465},
{-32'd6513, -32'd5407, 32'd3902, -32'd7428},
{-32'd1727, 32'd13427, -32'd6903, 32'd2006},
{-32'd5810, 32'd9265, 32'd8723, -32'd2634},
{32'd10127, 32'd508, 32'd492, 32'd2480},
{-32'd7345, 32'd121, -32'd5623, 32'd1787},
{-32'd11122, 32'd2886, -32'd9310, -32'd4181},
{-32'd9031, -32'd6973, -32'd2057, 32'd6244},
{32'd10449, 32'd2232, -32'd4491, 32'd8025},
{32'd2783, 32'd5411, 32'd8672, 32'd2380},
{32'd7677, 32'd2868, -32'd10532, 32'd3197},
{-32'd4677, -32'd2963, -32'd3347, -32'd922}
},
{{32'd1412, -32'd3931, 32'd7507, 32'd2820},
{32'd6449, -32'd12181, 32'd3695, 32'd3647},
{-32'd16769, -32'd2604, -32'd7563, -32'd487},
{32'd3194, 32'd3848, -32'd2994, 32'd7175},
{32'd7116, -32'd7139, 32'd2008, -32'd1933},
{-32'd7687, -32'd7585, -32'd4657, 32'd3487},
{32'd981, 32'd8267, 32'd5709, 32'd1314},
{-32'd3829, -32'd6817, 32'd1721, -32'd5826},
{32'd803, 32'd3471, -32'd35, 32'd16401},
{32'd14496, 32'd6635, 32'd1568, 32'd11497},
{32'd6748, -32'd2875, -32'd1710, -32'd2141},
{-32'd6839, 32'd7013, -32'd6190, -32'd7525},
{32'd2380, 32'd9723, -32'd12948, -32'd5021},
{32'd13060, 32'd4930, 32'd3091, -32'd8371},
{32'd9862, -32'd9858, 32'd4666, 32'd3330},
{32'd12767, -32'd7022, -32'd403, -32'd1126},
{-32'd2096, 32'd2098, 32'd13375, 32'd1035},
{32'd13018, 32'd16160, -32'd3449, -32'd2503},
{32'd8432, 32'd1491, 32'd149, 32'd2530},
{-32'd28, -32'd7078, 32'd8918, -32'd7882},
{-32'd7386, -32'd3654, -32'd868, 32'd3103},
{-32'd16323, -32'd13727, -32'd2032, -32'd5532},
{-32'd10943, -32'd5987, 32'd5738, 32'd4919},
{-32'd6426, -32'd5817, -32'd3214, -32'd9927},
{32'd3989, 32'd9225, -32'd4790, -32'd1301},
{-32'd6834, -32'd1986, -32'd6819, -32'd3942},
{-32'd12447, 32'd5006, 32'd6343, 32'd3335},
{32'd3054, -32'd8883, 32'd4156, -32'd1166},
{-32'd2746, 32'd2682, 32'd1579, -32'd825},
{-32'd7276, 32'd2765, -32'd5096, -32'd5383},
{32'd11442, -32'd10483, -32'd536, 32'd991},
{-32'd4099, -32'd10563, -32'd666, -32'd10892},
{32'd4514, 32'd1950, 32'd5384, 32'd8519},
{32'd6274, -32'd4688, -32'd12390, -32'd4158},
{32'd16111, 32'd7827, -32'd1551, 32'd12811},
{-32'd2577, -32'd8149, -32'd1050, -32'd11307},
{32'd9032, -32'd9467, -32'd5287, -32'd5107},
{32'd3944, -32'd4517, -32'd3521, 32'd854},
{-32'd3092, -32'd6333, 32'd5855, 32'd2293},
{32'd2393, -32'd4749, -32'd2186, -32'd627},
{-32'd2981, 32'd5701, 32'd5228, -32'd2314},
{-32'd1812, 32'd7212, -32'd2650, 32'd7810},
{-32'd1775, -32'd3121, 32'd3854, -32'd4655},
{32'd8305, -32'd2571, 32'd301, -32'd1913},
{-32'd5817, -32'd8835, -32'd5089, -32'd1401},
{32'd3784, 32'd1828, 32'd8559, 32'd8234},
{32'd5728, -32'd8917, -32'd10251, -32'd13228},
{32'd1500, 32'd3373, -32'd15494, -32'd7588},
{32'd7077, 32'd291, -32'd1698, -32'd6564},
{32'd1939, 32'd1126, -32'd354, -32'd8296},
{32'd1907, -32'd545, -32'd2081, 32'd2115},
{32'd8516, 32'd2385, -32'd9434, 32'd172},
{32'd7250, -32'd3091, 32'd2655, -32'd8145},
{-32'd3316, -32'd2644, 32'd2370, 32'd2573},
{-32'd1804, 32'd1376, 32'd6688, -32'd7740},
{32'd6630, -32'd10373, 32'd7797, -32'd269},
{32'd4887, -32'd3229, -32'd582, 32'd15542},
{32'd5128, -32'd14737, 32'd6161, -32'd5527},
{32'd7631, 32'd850, -32'd6246, -32'd11739},
{32'd1719, -32'd8335, 32'd198, -32'd3782},
{32'd1130, 32'd2864, -32'd4889, -32'd3578},
{-32'd3379, 32'd5827, 32'd1041, 32'd4231},
{32'd2943, -32'd8056, 32'd7044, -32'd14292},
{-32'd5045, 32'd592, 32'd7858, 32'd15060},
{-32'd4479, -32'd4983, -32'd6862, -32'd1953},
{-32'd3578, 32'd1216, 32'd97, 32'd5369},
{-32'd1494, 32'd3033, 32'd8287, 32'd4925},
{-32'd2815, -32'd9655, -32'd3797, -32'd6215},
{-32'd14925, 32'd13451, -32'd18, -32'd2739},
{32'd1530, -32'd7945, 32'd4796, 32'd12440},
{-32'd6042, -32'd8557, 32'd4513, 32'd4625},
{32'd5971, -32'd638, -32'd5475, -32'd7236},
{32'd4619, -32'd247, 32'd5447, 32'd2344},
{-32'd13793, 32'd2497, 32'd9340, 32'd1544},
{-32'd8413, 32'd6738, -32'd6050, 32'd2918},
{-32'd6355, 32'd17523, -32'd2894, 32'd4985},
{32'd6976, 32'd2445, -32'd4939, 32'd7421},
{-32'd9977, 32'd1605, 32'd4951, -32'd5138},
{-32'd1544, 32'd3170, -32'd11162, 32'd13},
{32'd3371, -32'd5032, 32'd1184, 32'd940},
{32'd1507, -32'd5762, -32'd934, -32'd1778},
{-32'd22729, 32'd3385, 32'd16182, 32'd1019},
{32'd22990, -32'd1425, -32'd6943, -32'd3160},
{-32'd7729, -32'd3701, 32'd1420, 32'd1392},
{32'd5408, 32'd4529, 32'd659, -32'd11987},
{-32'd4538, -32'd12464, 32'd15285, 32'd7121},
{-32'd6982, -32'd7277, -32'd6625, 32'd1391},
{32'd9298, -32'd1948, 32'd433, -32'd7519},
{-32'd4605, -32'd5079, -32'd10250, 32'd6473},
{-32'd1758, -32'd8751, -32'd2881, -32'd1831},
{32'd7453, 32'd4756, -32'd1800, 32'd3996},
{32'd2801, 32'd6531, 32'd3237, 32'd5900},
{32'd18656, -32'd253, -32'd4288, -32'd193},
{32'd12093, 32'd7885, -32'd1447, 32'd8856},
{-32'd9479, -32'd812, -32'd8993, 32'd1899},
{32'd405, -32'd12180, -32'd2930, 32'd14089},
{32'd4984, 32'd2459, 32'd3419, -32'd523},
{32'd13143, 32'd2974, -32'd6835, -32'd4823},
{32'd2532, -32'd1078, 32'd660, 32'd2655},
{32'd18865, -32'd1477, 32'd3290, -32'd1552},
{-32'd5158, -32'd12293, 32'd649, 32'd8645},
{-32'd16442, -32'd11841, 32'd5388, -32'd11934},
{32'd7230, -32'd3245, 32'd3387, 32'd1841},
{32'd10596, 32'd12639, 32'd709, -32'd418},
{-32'd12782, -32'd908, 32'd11734, 32'd6512},
{-32'd6955, -32'd4906, 32'd2369, 32'd10003},
{32'd1012, -32'd5314, 32'd716, 32'd1564},
{32'd1613, 32'd3557, 32'd4766, 32'd11226},
{32'd472, 32'd10967, -32'd645, -32'd3140},
{32'd865, -32'd1425, 32'd2037, 32'd3501},
{32'd832, -32'd67, -32'd1200, 32'd1988},
{-32'd5268, 32'd1007, 32'd7609, 32'd7652},
{32'd1895, 32'd1787, 32'd2032, -32'd1243},
{-32'd6497, 32'd6810, -32'd8583, -32'd4591},
{-32'd2681, -32'd4202, 32'd3403, -32'd11487},
{-32'd5361, -32'd2004, 32'd14399, 32'd5383},
{-32'd8758, 32'd6192, -32'd4763, -32'd6108},
{32'd629, -32'd9786, -32'd6962, -32'd319},
{32'd11512, -32'd5883, 32'd19427, -32'd6117},
{32'd12767, 32'd1845, 32'd7118, -32'd595},
{32'd4958, 32'd19808, 32'd914, 32'd129},
{-32'd2815, 32'd14954, -32'd4694, 32'd3774},
{-32'd6167, 32'd5173, 32'd11300, -32'd6011},
{-32'd17148, -32'd5910, 32'd2420, -32'd569},
{32'd1145, 32'd1392, -32'd6927, -32'd13838},
{-32'd7675, 32'd2678, 32'd602, -32'd1134},
{-32'd1916, 32'd4101, -32'd2098, -32'd1545},
{-32'd6126, -32'd8755, 32'd7132, 32'd2729},
{-32'd13256, -32'd4579, -32'd3462, -32'd445},
{32'd125, 32'd1152, -32'd2840, 32'd2929},
{-32'd8531, 32'd2038, 32'd10341, -32'd452},
{32'd2893, -32'd2382, -32'd5871, -32'd949},
{-32'd2232, -32'd2122, -32'd2388, 32'd2950},
{32'd4484, -32'd3456, 32'd5730, -32'd1285},
{-32'd6719, -32'd7362, -32'd8679, -32'd3912},
{-32'd10342, -32'd3632, 32'd3656, -32'd7302},
{-32'd4301, -32'd6711, -32'd12766, 32'd8984},
{-32'd7918, -32'd7285, -32'd10833, -32'd1871},
{-32'd1059, -32'd1551, 32'd7751, -32'd204},
{-32'd18676, -32'd7052, 32'd598, -32'd10055},
{-32'd15153, 32'd10863, -32'd5721, 32'd17462},
{-32'd8298, 32'd5236, -32'd3856, -32'd11674},
{32'd322, 32'd3658, 32'd7313, -32'd1084},
{-32'd7351, -32'd3901, -32'd1459, -32'd9834},
{32'd15351, 32'd2586, -32'd2405, -32'd2581},
{-32'd11467, 32'd3496, 32'd1908, 32'd6829},
{-32'd2585, -32'd418, -32'd4435, -32'd2896},
{32'd8203, -32'd2659, 32'd8645, -32'd1956},
{-32'd1162, 32'd8654, 32'd3702, 32'd4721},
{32'd3801, -32'd2417, -32'd1508, -32'd19174},
{32'd1798, -32'd5350, -32'd7669, -32'd10273},
{32'd4417, 32'd8808, 32'd10483, -32'd4058},
{32'd7423, 32'd5781, 32'd17444, -32'd675},
{32'd2996, -32'd3611, -32'd4062, 32'd7958},
{-32'd2382, -32'd9364, -32'd4818, -32'd11095},
{32'd4774, -32'd6616, 32'd5400, 32'd2718},
{32'd719, 32'd11183, -32'd4161, 32'd2291},
{32'd1199, 32'd7308, -32'd2299, 32'd3061},
{-32'd58, -32'd9336, 32'd4950, 32'd4009},
{-32'd7235, -32'd2875, -32'd7134, -32'd3638},
{-32'd3646, -32'd10155, 32'd1796, 32'd3860},
{32'd2361, 32'd5036, -32'd2586, 32'd10828},
{32'd120, -32'd4114, -32'd1342, -32'd7176},
{-32'd12100, 32'd2108, -32'd1316, 32'd4964},
{-32'd1228, 32'd6548, 32'd2788, 32'd3934},
{-32'd4635, -32'd3191, 32'd1116, -32'd5292},
{32'd10827, 32'd6056, -32'd5678, -32'd2419},
{-32'd6043, -32'd2961, -32'd216, -32'd262},
{-32'd6615, -32'd7789, -32'd4159, -32'd1063},
{-32'd3634, 32'd412, -32'd4002, 32'd2669},
{32'd1001, 32'd3063, -32'd5819, -32'd4678},
{-32'd2788, -32'd2326, -32'd7507, 32'd1619},
{32'd8768, 32'd4583, 32'd3912, 32'd12746},
{-32'd5739, -32'd8309, -32'd11658, -32'd1729},
{32'd4358, -32'd7681, -32'd1006, -32'd6756},
{32'd5413, -32'd2183, -32'd7832, 32'd1835},
{32'd2026, 32'd2342, 32'd4715, 32'd1090},
{-32'd5574, 32'd795, 32'd3680, 32'd5546},
{32'd1872, -32'd8237, 32'd15895, -32'd2489},
{-32'd14808, -32'd13724, -32'd3192, -32'd13167},
{-32'd26684, -32'd4478, 32'd10319, -32'd6809},
{32'd6193, -32'd5381, 32'd1283, 32'd1417},
{-32'd5164, -32'd5153, 32'd5711, -32'd12437},
{-32'd4297, -32'd161, -32'd12003, -32'd2451},
{-32'd2388, -32'd1788, -32'd6965, -32'd4459},
{-32'd4645, 32'd11299, -32'd5281, 32'd4056},
{-32'd4043, 32'd3054, -32'd3595, -32'd12829},
{-32'd2473, 32'd15747, 32'd10365, -32'd284},
{32'd8199, -32'd7589, -32'd277, 32'd24091},
{32'd5770, -32'd649, 32'd3555, -32'd10944},
{32'd653, 32'd7358, -32'd1746, -32'd8275},
{32'd7331, -32'd5331, 32'd7865, -32'd7250},
{32'd9936, 32'd1224, 32'd6408, 32'd8133},
{-32'd62, -32'd10222, 32'd906, -32'd1516},
{-32'd17496, 32'd4799, 32'd10409, 32'd5902},
{32'd10979, -32'd17904, 32'd6936, -32'd10549},
{-32'd7034, -32'd5902, -32'd1101, -32'd1653},
{32'd4411, -32'd3384, 32'd6040, 32'd2574},
{-32'd1437, -32'd7819, 32'd3902, -32'd7404},
{32'd9047, -32'd3142, -32'd292, 32'd10213},
{-32'd2516, -32'd10726, 32'd2289, -32'd11059},
{32'd2603, 32'd5372, -32'd2956, 32'd5657},
{-32'd4780, -32'd4986, 32'd3667, 32'd107},
{32'd2798, -32'd2976, 32'd10635, 32'd30},
{32'd4031, -32'd1590, -32'd7550, -32'd4774},
{32'd7537, 32'd926, -32'd431, -32'd6325},
{-32'd3406, -32'd1800, -32'd8394, 32'd17551},
{32'd20138, -32'd4174, -32'd5974, -32'd1860},
{-32'd2528, 32'd1211, -32'd8080, 32'd1955},
{-32'd5843, 32'd8818, -32'd6344, -32'd9179},
{-32'd4406, -32'd9554, -32'd10266, 32'd8654},
{-32'd13843, -32'd1995, 32'd6731, 32'd7087},
{-32'd18846, -32'd12650, -32'd2123, -32'd1927},
{32'd11346, 32'd13179, 32'd3401, 32'd5146},
{-32'd14875, -32'd8986, 32'd744, -32'd3323},
{32'd5209, -32'd3138, -32'd5811, 32'd1052},
{32'd1509, -32'd7375, -32'd9846, -32'd5228},
{-32'd7137, -32'd971, 32'd58, 32'd5543},
{-32'd7239, -32'd237, 32'd4920, -32'd6269},
{-32'd14404, -32'd7209, -32'd4046, 32'd2367},
{-32'd5987, -32'd1869, 32'd7395, -32'd2681},
{-32'd328, 32'd5848, 32'd1009, -32'd3620},
{-32'd6511, 32'd5745, -32'd1167, -32'd3118},
{-32'd9530, 32'd22360, 32'd6929, -32'd1310},
{32'd6375, -32'd7234, -32'd2484, -32'd2593},
{-32'd3598, -32'd4258, -32'd4276, 32'd4680},
{32'd437, -32'd570, -32'd6160, 32'd38},
{32'd3525, -32'd410, 32'd4840, 32'd6620},
{-32'd12312, 32'd6113, -32'd205, 32'd2099},
{32'd916, -32'd926, 32'd1063, 32'd5835},
{32'd3123, -32'd6468, 32'd56, 32'd5753},
{-32'd4717, -32'd2925, -32'd2554, -32'd823},
{32'd6827, -32'd3299, 32'd4447, -32'd4782},
{-32'd7195, -32'd5786, -32'd6696, 32'd5202},
{32'd11828, -32'd6076, -32'd87, -32'd8058},
{-32'd3586, -32'd10357, -32'd8554, -32'd5318},
{32'd9610, -32'd4855, 32'd2192, 32'd4999},
{32'd7115, -32'd3510, -32'd1379, -32'd2985},
{-32'd1243, 32'd9063, 32'd10074, -32'd1996},
{-32'd2433, 32'd8752, -32'd15620, -32'd3939},
{-32'd2039, -32'd2676, 32'd6422, -32'd258},
{-32'd4239, -32'd13313, -32'd6956, 32'd1606},
{32'd2598, -32'd6820, -32'd1368, -32'd5116},
{32'd1021, -32'd3760, -32'd9191, -32'd5814},
{32'd10418, 32'd15134, 32'd6768, 32'd9063},
{32'd15662, 32'd6543, 32'd2067, 32'd940},
{32'd8219, -32'd8214, -32'd857, -32'd9492},
{32'd8160, 32'd5047, -32'd14173, 32'd7227},
{32'd5880, -32'd3429, -32'd9069, 32'd1179},
{-32'd8759, -32'd17994, 32'd4273, 32'd8801},
{-32'd5335, 32'd6134, -32'd7577, 32'd10799},
{-32'd16353, 32'd11787, -32'd3972, 32'd2492},
{32'd4644, 32'd9558, 32'd9408, -32'd6794},
{32'd1657, -32'd9006, -32'd3716, 32'd6425},
{-32'd13955, 32'd2312, 32'd11557, 32'd7184},
{32'd856, -32'd1870, 32'd3319, 32'd1825},
{32'd9756, 32'd4786, 32'd1478, 32'd4464},
{32'd4406, 32'd2586, 32'd2611, 32'd8179},
{32'd1181, 32'd3925, 32'd381, -32'd707},
{32'd1503, 32'd5728, 32'd2456, -32'd476},
{32'd7199, -32'd8089, -32'd1248, -32'd4524},
{32'd13596, 32'd7154, -32'd5455, -32'd3617},
{-32'd23137, -32'd15386, 32'd5059, -32'd3275},
{-32'd12729, 32'd262, -32'd7430, -32'd2120},
{32'd806, 32'd1471, 32'd876, 32'd8128},
{-32'd20237, -32'd6626, 32'd3399, 32'd6260},
{32'd7920, 32'd8013, -32'd5409, 32'd421},
{32'd9685, 32'd4945, -32'd4844, -32'd2066},
{-32'd861, -32'd1218, -32'd995, -32'd18614},
{32'd4607, -32'd3419, 32'd3225, 32'd1790},
{32'd5942, 32'd258, 32'd1300, -32'd101},
{32'd423, 32'd3400, -32'd3631, 32'd6383},
{-32'd1295, -32'd5377, 32'd5215, -32'd1790},
{32'd5605, 32'd5481, 32'd2155, -32'd1183},
{-32'd1056, 32'd1067, 32'd1491, -32'd4495},
{32'd10066, 32'd591, 32'd2623, 32'd2018},
{32'd17159, 32'd10228, 32'd1083, 32'd11670},
{32'd1419, 32'd12746, 32'd10684, -32'd9514},
{-32'd7256, -32'd7114, 32'd2887, -32'd2662},
{32'd5276, 32'd3307, -32'd5066, 32'd2451},
{-32'd1102, 32'd2307, -32'd1883, 32'd10908},
{-32'd9676, 32'd5842, 32'd9585, 32'd5177},
{-32'd8670, 32'd9813, 32'd12534, 32'd11759},
{-32'd5347, -32'd7329, -32'd6304, 32'd1564},
{32'd5219, -32'd2478, 32'd1615, 32'd1803},
{-32'd991, -32'd5688, -32'd5084, -32'd8980},
{32'd3584, 32'd6475, 32'd13681, 32'd7171},
{-32'd9934, 32'd1207, 32'd10282, -32'd5256},
{32'd11755, 32'd5887, -32'd4113, 32'd799},
{32'd10512, -32'd4885, 32'd8617, 32'd1100},
{-32'd4413, -32'd644, -32'd5725, 32'd2655},
{32'd1342, 32'd3443, -32'd7394, -32'd1070},
{-32'd396, -32'd4589, 32'd2032, 32'd5951},
{-32'd9057, 32'd3065, 32'd1087, -32'd111},
{32'd2348, 32'd1819, 32'd13165, -32'd2083},
{-32'd1538, 32'd1107, -32'd7320, -32'd5065},
{32'd12622, 32'd20, -32'd4518, 32'd15848},
{32'd6572, -32'd216, 32'd1307, 32'd3785},
{32'd5416, -32'd1689, -32'd4578, -32'd4142},
{32'd6611, 32'd11199, -32'd406, -32'd1312}
},
{{-32'd1368, 32'd4048, -32'd4460, -32'd674},
{32'd7507, 32'd2416, 32'd4242, 32'd8124},
{-32'd11866, 32'd13450, -32'd5065, -32'd7236},
{32'd6968, -32'd4195, -32'd16126, 32'd7029},
{-32'd2575, 32'd6958, 32'd2299, 32'd1127},
{-32'd4648, -32'd1990, -32'd1950, 32'd1089},
{32'd1594, 32'd13156, 32'd5251, 32'd8282},
{32'd436, -32'd444, -32'd5282, 32'd353},
{32'd12227, 32'd8603, 32'd3199, -32'd9203},
{-32'd1283, 32'd25, -32'd1489, 32'd6316},
{32'd5840, 32'd3398, -32'd4282, -32'd3269},
{-32'd9933, -32'd1106, -32'd6087, 32'd8602},
{-32'd286, 32'd9309, -32'd9696, 32'd3966},
{-32'd4622, -32'd2736, -32'd10451, -32'd1641},
{-32'd181, -32'd2428, 32'd2598, 32'd4108},
{32'd782, -32'd1337, 32'd4663, -32'd10889},
{32'd7525, 32'd1732, -32'd4217, 32'd9494},
{-32'd5778, 32'd7778, 32'd13538, 32'd8774},
{-32'd12721, -32'd22384, -32'd15838, -32'd10609},
{-32'd5547, -32'd4354, -32'd1309, 32'd4036},
{-32'd8182, 32'd1588, -32'd6415, -32'd3323},
{-32'd14282, -32'd6684, -32'd9208, 32'd7361},
{-32'd4629, -32'd5360, 32'd41, 32'd1919},
{32'd2409, 32'd134, -32'd1503, -32'd16895},
{32'd6565, 32'd8007, -32'd3364, 32'd2490},
{32'd1280, 32'd2403, -32'd4372, 32'd4867},
{32'd641, 32'd260, -32'd9384, -32'd5108},
{-32'd2053, 32'd14844, 32'd8224, -32'd5850},
{32'd1262, 32'd811, -32'd4807, 32'd2900},
{-32'd16692, -32'd8770, -32'd9113, -32'd5517},
{-32'd12718, -32'd13238, -32'd10054, 32'd2253},
{-32'd6405, -32'd11917, 32'd846, -32'd5680},
{-32'd4638, 32'd2665, 32'd5220, 32'd6892},
{-32'd3634, -32'd4068, 32'd2522, -32'd3505},
{-32'd3531, 32'd6419, 32'd522, 32'd5382},
{32'd5055, 32'd3499, 32'd7958, -32'd398},
{-32'd4740, 32'd7553, 32'd682, 32'd8262},
{-32'd5942, 32'd7286, 32'd12186, -32'd234},
{32'd13976, 32'd7908, 32'd1646, -32'd7927},
{32'd5618, 32'd3794, 32'd8113, 32'd293},
{-32'd2354, 32'd5821, 32'd1595, 32'd12114},
{-32'd3084, 32'd4970, 32'd6631, -32'd470},
{32'd4696, -32'd107, 32'd20515, -32'd1711},
{-32'd3778, -32'd4106, 32'd6188, -32'd9541},
{32'd1853, 32'd3406, -32'd3839, 32'd819},
{32'd4946, 32'd3966, -32'd2191, -32'd2900},
{-32'd16269, -32'd4548, -32'd1352, -32'd5317},
{-32'd11865, -32'd12408, -32'd6506, -32'd5218},
{32'd7824, 32'd12089, -32'd9719, 32'd3119},
{-32'd10218, 32'd1074, 32'd18719, 32'd14501},
{32'd5724, -32'd10000, -32'd10822, 32'd6981},
{32'd5115, 32'd5722, 32'd15045, 32'd2743},
{-32'd8744, 32'd6226, -32'd13756, -32'd5498},
{-32'd9374, 32'd6196, 32'd5158, 32'd1839},
{32'd6237, 32'd7522, -32'd7888, 32'd6201},
{32'd6107, 32'd6141, 32'd2920, 32'd12792},
{-32'd4632, 32'd2420, -32'd5577, -32'd1310},
{32'd274, -32'd8843, -32'd500, 32'd2786},
{32'd3008, 32'd1534, 32'd8934, -32'd923},
{-32'd6138, 32'd7715, -32'd489, 32'd1369},
{32'd59, 32'd2094, -32'd19122, 32'd2122},
{32'd12416, 32'd11382, 32'd4088, -32'd14815},
{32'd301, -32'd3016, -32'd3037, 32'd845},
{-32'd6139, -32'd5940, 32'd2584, -32'd5231},
{-32'd6478, 32'd1018, 32'd567, -32'd4531},
{32'd12810, 32'd7004, -32'd877, 32'd3770},
{-32'd6238, -32'd9461, -32'd13119, -32'd4699},
{-32'd2917, 32'd318, 32'd938, -32'd8552},
{32'd2979, -32'd561, -32'd14674, -32'd2238},
{-32'd909, 32'd2385, -32'd2741, 32'd6123},
{-32'd2261, 32'd9804, 32'd6222, -32'd2675},
{-32'd831, 32'd2322, 32'd9874, -32'd218},
{32'd9911, -32'd3265, -32'd5273, -32'd4739},
{-32'd2719, -32'd8435, 32'd5928, 32'd3673},
{32'd1648, -32'd2546, -32'd10742, 32'd7590},
{32'd757, 32'd11441, 32'd17075, -32'd12327},
{-32'd7144, -32'd6407, 32'd10403, -32'd7063},
{-32'd10740, -32'd6155, -32'd7545, -32'd10136},
{32'd5094, 32'd1411, -32'd6075, 32'd28},
{-32'd3364, 32'd3696, -32'd6395, -32'd1400},
{-32'd820, 32'd6867, -32'd3869, -32'd6755},
{32'd6589, 32'd935, 32'd3752, -32'd2537},
{32'd4631, -32'd1884, -32'd2980, 32'd1780},
{-32'd235, 32'd2902, 32'd10874, 32'd7900},
{-32'd9854, -32'd2436, 32'd2644, 32'd626},
{-32'd5820, -32'd4376, -32'd14208, 32'd284},
{-32'd16373, 32'd2842, -32'd5810, -32'd4453},
{-32'd7391, -32'd3914, -32'd1770, -32'd11580},
{32'd11627, 32'd2095, -32'd10310, -32'd4040},
{-32'd818, -32'd4167, -32'd15426, 32'd998},
{32'd1467, 32'd5427, 32'd6399, 32'd10251},
{32'd1693, 32'd4418, 32'd6357, 32'd3434},
{32'd9017, 32'd11931, 32'd1014, -32'd10627},
{-32'd14399, 32'd10957, -32'd4546, -32'd1899},
{32'd12031, 32'd8243, 32'd7096, 32'd4511},
{32'd856, 32'd10853, 32'd1299, 32'd1946},
{-32'd421, 32'd1221, 32'd4387, 32'd2869},
{-32'd4641, 32'd5922, 32'd7813, 32'd5272},
{-32'd4288, 32'd15734, 32'd5667, -32'd4676},
{-32'd982, 32'd1298, 32'd11445, 32'd2809},
{-32'd10154, -32'd11862, 32'd19619, -32'd3789},
{-32'd6659, -32'd5539, 32'd9510, 32'd2268},
{32'd4757, 32'd5044, -32'd2794, -32'd4685},
{32'd1878, -32'd3179, 32'd2368, -32'd13822},
{-32'd4666, -32'd1061, 32'd23646, 32'd12397},
{-32'd4542, 32'd476, 32'd827, -32'd3146},
{-32'd9349, -32'd6, -32'd3360, -32'd2213},
{-32'd9035, 32'd1365, -32'd2265, -32'd6795},
{-32'd5400, -32'd6461, -32'd14191, 32'd6248},
{-32'd18282, -32'd1201, 32'd2091, 32'd141},
{32'd13475, 32'd25798, -32'd6126, 32'd2068},
{32'd6640, 32'd3848, 32'd3625, -32'd4748},
{32'd3614, 32'd9136, -32'd5900, 32'd4430},
{-32'd681, 32'd1897, -32'd3060, 32'd6557},
{32'd1642, -32'd7884, -32'd4366, 32'd1285},
{32'd7971, 32'd1527, 32'd13487, 32'd1503},
{-32'd5263, 32'd11098, 32'd10616, 32'd14972},
{32'd1406, 32'd10097, 32'd17765, 32'd6034},
{-32'd4555, 32'd5860, 32'd13156, -32'd3959},
{32'd10119, 32'd4551, 32'd1843, 32'd3086},
{-32'd290, 32'd6088, -32'd8024, -32'd4805},
{32'd6173, 32'd7188, -32'd1790, -32'd3494},
{32'd6026, 32'd8606, 32'd4691, 32'd10093},
{32'd6444, 32'd3232, 32'd11262, 32'd5819},
{-32'd21598, -32'd5500, -32'd9111, -32'd3991},
{32'd7447, 32'd3876, -32'd7469, 32'd399},
{32'd17589, -32'd5302, -32'd7038, 32'd13358},
{-32'd3911, 32'd12006, -32'd1240, -32'd3989},
{-32'd10308, -32'd6948, 32'd2719, 32'd6620},
{32'd2618, 32'd10816, 32'd1914, 32'd3123},
{-32'd3665, -32'd2374, 32'd7964, 32'd9310},
{32'd6346, 32'd1421, 32'd9608, 32'd978},
{-32'd1640, 32'd1754, -32'd2204, -32'd7717},
{32'd16523, 32'd6930, 32'd10543, -32'd4010},
{-32'd3610, -32'd2729, -32'd241, -32'd2579},
{32'd4324, 32'd4493, -32'd1881, 32'd2329},
{32'd8640, 32'd256, -32'd208, 32'd2901},
{32'd4475, 32'd855, 32'd9917, 32'd3633},
{32'd4883, 32'd327, -32'd6479, -32'd2787},
{-32'd3634, -32'd4972, 32'd13976, 32'd10461},
{-32'd4888, 32'd2505, 32'd9604, -32'd10675},
{32'd7124, 32'd3297, 32'd5544, -32'd9282},
{32'd11320, -32'd94, -32'd2131, -32'd509},
{-32'd13170, -32'd1631, 32'd6111, 32'd3091},
{-32'd929, 32'd7226, -32'd4478, -32'd1480},
{32'd14359, 32'd10853, 32'd17667, 32'd9420},
{-32'd4532, -32'd10001, 32'd7642, -32'd11544},
{-32'd5395, -32'd2787, -32'd202, 32'd5441},
{32'd11409, 32'd3714, 32'd11539, 32'd9841},
{-32'd11333, -32'd9601, -32'd2085, 32'd2397},
{-32'd1717, 32'd129, 32'd3329, -32'd7600},
{32'd10768, -32'd8795, 32'd1234, 32'd2551},
{-32'd3755, -32'd5935, 32'd1389, 32'd11077},
{-32'd718, 32'd6436, -32'd6148, 32'd3339},
{-32'd14317, 32'd1761, 32'd567, -32'd10377},
{-32'd1622, -32'd10543, 32'd958, -32'd1213},
{-32'd7176, -32'd11601, -32'd998, -32'd1797},
{-32'd4577, -32'd3891, -32'd15488, 32'd7223},
{-32'd8508, -32'd10785, -32'd8835, -32'd4842},
{-32'd2722, 32'd763, 32'd2160, 32'd5432},
{-32'd472, -32'd4338, 32'd256, -32'd8064},
{32'd2908, -32'd2606, 32'd2433, 32'd1964},
{-32'd2137, -32'd2841, 32'd2620, -32'd1005},
{32'd6545, 32'd9201, -32'd449, -32'd323},
{-32'd59, 32'd10557, 32'd17140, 32'd12159},
{-32'd4757, -32'd6802, -32'd1575, 32'd11042},
{-32'd8284, 32'd664, 32'd8825, 32'd3564},
{32'd5022, 32'd4151, -32'd1374, 32'd5760},
{32'd1646, 32'd1418, 32'd7345, 32'd996},
{-32'd17231, -32'd6701, 32'd475, -32'd56},
{-32'd6594, 32'd2682, 32'd1519, 32'd4200},
{-32'd4531, -32'd2876, 32'd5894, 32'd4341},
{32'd4011, 32'd4513, -32'd741, -32'd1900},
{32'd1741, -32'd6913, -32'd6543, -32'd9565},
{32'd4077, 32'd3542, -32'd11159, 32'd6490},
{-32'd19303, -32'd6249, -32'd5765, 32'd6110},
{32'd20825, -32'd4833, 32'd4662, 32'd1289},
{-32'd130, 32'd3283, -32'd4243, -32'd7952},
{-32'd2203, -32'd5300, 32'd14698, -32'd242},
{-32'd12295, -32'd766, -32'd5769, -32'd2847},
{32'd4008, 32'd4010, 32'd4934, -32'd2122},
{-32'd6521, -32'd10663, 32'd7002, -32'd13510},
{-32'd3448, -32'd4269, 32'd4828, -32'd16282},
{32'd11854, 32'd2149, -32'd2887, -32'd3163},
{-32'd5995, 32'd9991, -32'd885, -32'd2091},
{32'd885, -32'd45, -32'd7933, 32'd4824},
{32'd9009, 32'd4142, 32'd10816, 32'd12481},
{32'd6605, -32'd5730, 32'd18058, -32'd7822},
{32'd6320, 32'd477, 32'd8925, -32'd15838},
{-32'd4391, -32'd3440, -32'd7985, 32'd1044},
{-32'd3844, 32'd3115, 32'd20813, 32'd340},
{32'd8233, -32'd4845, 32'd6987, -32'd1550},
{32'd1996, 32'd5220, -32'd6518, -32'd16606},
{-32'd1771, 32'd1384, -32'd5264, -32'd2897},
{32'd1869, -32'd7888, -32'd1710, -32'd11615},
{-32'd455, -32'd16532, -32'd7809, 32'd4512},
{-32'd3356, -32'd8308, 32'd13193, -32'd4008},
{32'd12983, 32'd3478, 32'd5186, -32'd37},
{32'd2596, -32'd1822, -32'd3736, -32'd6520},
{32'd8788, 32'd7916, 32'd12406, 32'd2359},
{-32'd8551, -32'd6928, -32'd2492, -32'd6384},
{-32'd2115, 32'd18254, -32'd5612, 32'd1594},
{-32'd593, -32'd2226, 32'd6036, -32'd1213},
{32'd11081, -32'd9251, -32'd7311, 32'd8446},
{32'd2769, -32'd5696, 32'd1855, -32'd4200},
{-32'd5296, 32'd3997, -32'd4186, 32'd985},
{32'd13979, -32'd1021, 32'd9375, -32'd143},
{32'd2611, 32'd6875, -32'd6307, 32'd1456},
{-32'd8658, 32'd3388, -32'd17091, -32'd1005},
{32'd11685, 32'd3475, 32'd5671, -32'd2880},
{-32'd745, 32'd12953, -32'd7795, -32'd2774},
{-32'd8224, 32'd5683, 32'd2758, 32'd4810},
{-32'd3794, -32'd4516, -32'd3936, 32'd5304},
{32'd7457, 32'd10194, 32'd3226, -32'd713},
{-32'd1057, -32'd8985, -32'd10692, -32'd6984},
{-32'd21269, -32'd9405, -32'd7960, -32'd1994},
{32'd6809, 32'd6910, 32'd240, -32'd4774},
{32'd2421, -32'd8418, -32'd10681, -32'd823},
{32'd7666, 32'd4675, 32'd8017, 32'd15990},
{32'd2619, 32'd652, -32'd6070, -32'd2134},
{-32'd7284, 32'd2619, 32'd6109, -32'd3501},
{32'd6287, -32'd3368, 32'd11374, -32'd5499},
{-32'd1544, -32'd5152, -32'd4754, -32'd9650},
{32'd11162, -32'd7099, -32'd7238, 32'd9932},
{-32'd1604, -32'd2859, -32'd18758, -32'd3235},
{32'd6221, -32'd10482, -32'd7391, 32'd212},
{-32'd3705, -32'd4357, 32'd971, -32'd6162},
{32'd10942, -32'd1793, -32'd4770, -32'd7169},
{-32'd4338, -32'd3900, 32'd7249, 32'd2742},
{32'd5505, 32'd9737, -32'd4521, 32'd9652},
{-32'd9031, -32'd7432, -32'd445, 32'd2156},
{32'd1497, 32'd2189, -32'd791, 32'd4215},
{-32'd10700, -32'd3984, -32'd9676, -32'd3928},
{-32'd3222, 32'd90, -32'd8051, -32'd2953},
{32'd740, 32'd2667, 32'd8980, 32'd2259},
{32'd4775, -32'd4880, -32'd5114, -32'd2580},
{-32'd6663, 32'd3305, 32'd934, 32'd8082},
{32'd281, -32'd2807, -32'd1928, -32'd2974},
{32'd3455, 32'd6426, 32'd1531, -32'd12913},
{32'd1247, 32'd16132, -32'd2326, 32'd4951},
{32'd6941, 32'd3916, 32'd11728, -32'd1594},
{32'd3982, 32'd592, -32'd11019, -32'd922},
{-32'd895, 32'd3500, -32'd3541, -32'd1913},
{32'd5506, 32'd6507, 32'd1358, 32'd31},
{-32'd3198, -32'd4855, -32'd890, -32'd661},
{32'd1820, -32'd7019, -32'd878, -32'd10088},
{-32'd5596, 32'd553, 32'd11642, -32'd3033},
{-32'd4357, -32'd5718, -32'd7988, -32'd6248},
{-32'd14626, -32'd12619, -32'd6687, -32'd2646},
{-32'd3688, -32'd6982, -32'd2823, 32'd1266},
{-32'd9067, -32'd994, 32'd244, -32'd2734},
{-32'd11333, -32'd5949, -32'd10074, 32'd6271},
{32'd7771, 32'd2596, 32'd6842, 32'd1936},
{32'd65, -32'd8138, -32'd12974, -32'd6089},
{32'd3948, -32'd4966, 32'd9712, -32'd1901},
{32'd3030, -32'd10448, 32'd2360, 32'd4094},
{32'd254, -32'd6199, -32'd13392, -32'd13691},
{32'd12024, -32'd887, -32'd14697, 32'd179},
{32'd12051, -32'd2552, 32'd12322, 32'd3887},
{32'd9302, 32'd15618, 32'd4406, -32'd3029},
{-32'd10024, -32'd4229, -32'd20816, 32'd13423},
{-32'd5046, -32'd2740, -32'd10327, -32'd5288},
{-32'd8629, -32'd6145, 32'd6814, -32'd12484},
{32'd2501, 32'd17308, 32'd4345, -32'd5809},
{32'd4400, 32'd10677, 32'd3852, -32'd878},
{32'd3996, 32'd3022, -32'd7542, -32'd2391},
{32'd7803, -32'd8564, -32'd4952, 32'd6605},
{-32'd8321, 32'd1662, -32'd7302, 32'd7352},
{-32'd1938, 32'd10291, 32'd5426, -32'd282},
{32'd3607, -32'd7924, 32'd3663, -32'd2994},
{32'd2080, 32'd9818, -32'd2138, -32'd2117},
{32'd1997, -32'd678, -32'd7851, 32'd2030},
{-32'd15060, -32'd8571, -32'd1931, -32'd4485},
{32'd5998, 32'd4280, 32'd16816, -32'd1967},
{32'd3679, 32'd1779, 32'd7038, -32'd1979},
{-32'd6544, 32'd1674, -32'd7928, -32'd8046},
{-32'd2441, 32'd2077, -32'd1225, 32'd7367},
{32'd2318, 32'd12207, 32'd3630, 32'd5045},
{32'd1291, -32'd10584, -32'd6038, -32'd6823},
{-32'd4076, -32'd9441, 32'd4166, 32'd1310},
{-32'd989, -32'd386, -32'd8129, -32'd10615},
{32'd228, 32'd10875, 32'd12952, 32'd2962},
{32'd1216, -32'd3747, 32'd5868, -32'd702},
{-32'd240, 32'd862, 32'd4919, -32'd61},
{32'd5948, 32'd11635, -32'd8335, 32'd789},
{32'd819, -32'd3358, -32'd5656, 32'd2996},
{32'd6088, 32'd619, -32'd5292, 32'd10197},
{-32'd8612, -32'd11557, -32'd11279, -32'd4973},
{-32'd1798, 32'd4539, 32'd20171, -32'd5908},
{32'd3517, -32'd9112, 32'd10207, 32'd6102},
{-32'd12789, -32'd9448, -32'd8082, -32'd961},
{32'd707, 32'd5472, 32'd1780, 32'd3732},
{32'd11144, -32'd4071, -32'd8235, -32'd5569},
{-32'd937, -32'd9891, 32'd2203, -32'd7891},
{32'd4741, -32'd3024, 32'd5096, 32'd2636},
{-32'd2553, 32'd2532, 32'd1274, 32'd880},
{32'd9135, -32'd1526, -32'd2684, -32'd2898},
{32'd1177, 32'd1350, -32'd925, 32'd10906},
{32'd1396, -32'd579, -32'd14128, -32'd1893},
{32'd96, -32'd8278, 32'd6238, -32'd2594}
},
{{32'd8331, 32'd3198, 32'd944, -32'd179},
{-32'd3326, -32'd4282, -32'd8015, 32'd1997},
{-32'd8495, -32'd17488, -32'd2128, -32'd2397},
{32'd13551, 32'd5582, -32'd2836, 32'd1412},
{-32'd2657, 32'd2389, 32'd2922, 32'd968},
{-32'd140, 32'd10219, -32'd14000, 32'd16706},
{32'd595, -32'd226, -32'd5859, 32'd3438},
{32'd11816, 32'd3586, -32'd15504, -32'd3394},
{32'd10943, 32'd1753, 32'd18160, 32'd8205},
{32'd11967, 32'd5814, 32'd283, 32'd1290},
{-32'd5226, -32'd2101, -32'd1338, 32'd3507},
{32'd7110, -32'd6617, 32'd8994, -32'd5385},
{-32'd1096, 32'd696, 32'd6271, 32'd6326},
{-32'd3506, 32'd407, -32'd8524, -32'd5399},
{-32'd9457, -32'd3431, -32'd7646, -32'd888},
{-32'd8903, -32'd5335, 32'd4823, -32'd906},
{32'd3374, 32'd8767, 32'd1299, 32'd3240},
{32'd3636, -32'd6303, 32'd4123, -32'd8696},
{32'd7346, -32'd2053, -32'd13220, -32'd1297},
{32'd5229, -32'd5403, -32'd1769, 32'd8981},
{-32'd3826, 32'd2501, -32'd11435, 32'd5297},
{-32'd5283, 32'd505, -32'd4027, 32'd4364},
{-32'd14848, 32'd6133, -32'd1768, 32'd4346},
{-32'd8633, -32'd2580, 32'd7184, -32'd3152},
{32'd3570, -32'd829, -32'd6978, 32'd2622},
{-32'd1523, -32'd13079, -32'd9467, 32'd5186},
{-32'd3504, -32'd1384, 32'd4409, -32'd1133},
{-32'd6922, 32'd8923, 32'd1244, -32'd2839},
{-32'd2709, -32'd326, 32'd1129, 32'd2516},
{32'd3832, -32'd8294, -32'd523, -32'd1335},
{-32'd3066, -32'd7660, 32'd1570, 32'd10030},
{32'd3768, -32'd1935, -32'd1840, 32'd3415},
{32'd5142, 32'd6463, 32'd5568, -32'd4848},
{-32'd2152, -32'd4452, 32'd1613, -32'd5768},
{32'd2142, 32'd4604, -32'd773, 32'd2853},
{-32'd826, -32'd5001, -32'd2722, -32'd2416},
{-32'd283, 32'd10386, 32'd7012, -32'd13246},
{32'd2398, -32'd6138, 32'd8601, 32'd725},
{32'd7570, -32'd8807, 32'd8289, 32'd158},
{-32'd5293, 32'd1745, -32'd2921, 32'd5501},
{-32'd5424, 32'd538, 32'd7353, -32'd5593},
{32'd4957, -32'd3425, 32'd2485, 32'd1860},
{32'd778, -32'd1736, 32'd7233, -32'd13803},
{-32'd5314, -32'd5106, -32'd4388, -32'd878},
{-32'd2023, -32'd4085, 32'd1104, 32'd529},
{32'd2479, -32'd155, 32'd2509, 32'd2983},
{-32'd1686, -32'd10090, -32'd8893, -32'd343},
{-32'd4288, -32'd12108, 32'd5614, -32'd5973},
{32'd2553, 32'd9334, 32'd1253, -32'd2737},
{32'd1787, -32'd10244, -32'd5906, -32'd8415},
{32'd501, 32'd7208, 32'd18305, -32'd2346},
{32'd1361, 32'd4561, 32'd3948, -32'd9492},
{-32'd15127, -32'd2808, -32'd1793, -32'd5857},
{-32'd4170, -32'd8539, 32'd2117, -32'd5778},
{32'd9317, 32'd5241, 32'd2828, -32'd2994},
{32'd2461, 32'd221, -32'd9191, 32'd4925},
{32'd4456, -32'd7864, 32'd7930, -32'd1567},
{32'd4456, -32'd4655, 32'd3227, -32'd9241},
{-32'd16906, -32'd6173, 32'd4879, -32'd3460},
{32'd183, -32'd1157, 32'd2209, 32'd8680},
{-32'd270, -32'd1660, -32'd4291, 32'd5222},
{-32'd2088, 32'd12528, 32'd2667, 32'd1395},
{-32'd4294, 32'd1496, 32'd680, -32'd1451},
{32'd1898, 32'd1157, -32'd8186, 32'd6950},
{32'd1861, -32'd3789, -32'd2431, -32'd3570},
{-32'd240, -32'd4995, -32'd1915, 32'd87},
{32'd308, -32'd1799, 32'd2878, 32'd3327},
{-32'd6449, -32'd6538, 32'd1542, 32'd1663},
{-32'd146, -32'd14053, -32'd3905, 32'd1489},
{-32'd7529, 32'd10541, -32'd873, -32'd1071},
{-32'd4501, 32'd3472, 32'd69, 32'd1631},
{-32'd9425, 32'd1684, -32'd2796, -32'd7835},
{-32'd951, -32'd8039, -32'd1298, -32'd1723},
{-32'd2229, 32'd1411, -32'd5697, 32'd13051},
{32'd1703, 32'd978, 32'd136, 32'd10308},
{32'd6622, -32'd660, 32'd8308, -32'd4135},
{-32'd1188, -32'd4161, -32'd830, -32'd7009},
{32'd2300, 32'd358, 32'd6164, 32'd2541},
{32'd1345, -32'd614, 32'd7110, 32'd182},
{32'd3711, -32'd1054, -32'd99, -32'd7985},
{-32'd464, 32'd4933, 32'd3487, -32'd10286},
{32'd5376, -32'd5145, -32'd7674, -32'd4348},
{-32'd3200, 32'd2077, -32'd4373, 32'd3507},
{32'd8072, 32'd1631, 32'd14093, -32'd1509},
{32'd759, -32'd21025, 32'd2651, -32'd4776},
{-32'd6545, 32'd397, -32'd9669, -32'd4525},
{32'd1324, -32'd717, 32'd4220, -32'd5598},
{-32'd7800, -32'd1528, 32'd1294, -32'd4237},
{32'd4093, -32'd11710, 32'd10689, 32'd2557},
{32'd2131, -32'd1920, -32'd2298, -32'd2113},
{32'd6841, 32'd7279, 32'd256, -32'd1183},
{-32'd8385, -32'd3412, -32'd8372, 32'd10321},
{-32'd9437, -32'd6048, -32'd11183, 32'd383},
{-32'd5029, -32'd1790, 32'd8949, 32'd4292},
{-32'd831, 32'd1184, -32'd3792, 32'd4892},
{32'd1854, -32'd11816, 32'd1434, 32'd286},
{32'd1364, 32'd4611, 32'd987, -32'd241},
{-32'd1565, 32'd2878, -32'd3590, 32'd240},
{-32'd11570, -32'd686, 32'd6238, 32'd13579},
{32'd5039, 32'd7988, 32'd880, 32'd1040},
{-32'd15128, -32'd3047, -32'd15041, -32'd1819},
{-32'd4073, -32'd920, 32'd2959, 32'd2664},
{-32'd17039, 32'd14606, -32'd2214, 32'd1072},
{32'd2188, -32'd1950, 32'd4275, 32'd3602},
{-32'd4752, 32'd9266, 32'd7145, 32'd440},
{-32'd961, 32'd974, -32'd8165, -32'd1416},
{-32'd9301, 32'd6383, -32'd6099, 32'd1902},
{-32'd10036, -32'd265, 32'd2627, 32'd4714},
{-32'd2414, 32'd8855, 32'd6623, 32'd3567},
{32'd3809, -32'd6739, -32'd2191, 32'd3031},
{-32'd2453, -32'd5178, 32'd8089, -32'd7905},
{32'd1408, 32'd12069, 32'd1782, 32'd791},
{-32'd2535, -32'd4486, 32'd5975, 32'd1772},
{-32'd1668, 32'd3264, 32'd1934, 32'd11381},
{32'd2607, -32'd4112, -32'd2336, 32'd1279},
{32'd464, 32'd5328, -32'd602, 32'd367},
{-32'd3431, 32'd322, 32'd1511, 32'd773},
{-32'd609, 32'd4907, -32'd2772, 32'd4449},
{32'd1494, 32'd8967, -32'd1260, -32'd15327},
{32'd1670, 32'd4421, 32'd59, -32'd4663},
{-32'd6221, -32'd11129, -32'd9486, -32'd2740},
{-32'd3655, -32'd876, 32'd4522, -32'd5752},
{32'd2739, 32'd3439, -32'd2524, 32'd6707},
{-32'd959, -32'd11392, 32'd5398, 32'd11881},
{-32'd1134, -32'd4867, -32'd3566, -32'd9},
{-32'd4259, 32'd604, -32'd2288, 32'd4655},
{32'd7663, 32'd1746, -32'd10696, 32'd6722},
{-32'd4613, -32'd3401, -32'd6319, -32'd2761},
{32'd6058, 32'd591, -32'd4978, 32'd8767},
{-32'd8171, -32'd11975, 32'd5283, 32'd2725},
{-32'd2449, -32'd1889, -32'd5512, -32'd1662},
{32'd1634, -32'd4905, 32'd660, 32'd8296},
{-32'd6593, -32'd2580, -32'd1608, -32'd1451},
{32'd9086, 32'd7298, -32'd7692, 32'd9954},
{-32'd2319, -32'd1421, 32'd1656, -32'd3086},
{-32'd4985, -32'd4816, -32'd5102, 32'd1150},
{32'd1617, -32'd2685, 32'd3123, 32'd546},
{32'd375, -32'd11715, 32'd7993, -32'd216},
{32'd4196, -32'd1182, 32'd5199, 32'd3694},
{-32'd14814, 32'd741, -32'd3372, -32'd25},
{-32'd2795, 32'd1154, 32'd441, -32'd2134},
{-32'd7991, -32'd3162, 32'd1541, 32'd2212},
{32'd4054, 32'd6459, -32'd9818, -32'd9628},
{32'd1079, -32'd5474, 32'd3954, 32'd356},
{32'd8423, -32'd1830, 32'd1586, -32'd3362},
{32'd2072, 32'd11523, -32'd2058, -32'd8080},
{-32'd7112, -32'd423, -32'd8801, 32'd3956},
{-32'd2186, -32'd7395, -32'd16210, 32'd11883},
{32'd11471, -32'd224, -32'd1071, 32'd1969},
{-32'd5223, 32'd175, -32'd9505, -32'd5389},
{-32'd9209, 32'd1369, 32'd5504, -32'd9684},
{32'd293, 32'd16380, -32'd2099, -32'd12807},
{-32'd8865, 32'd4412, 32'd12, -32'd1290},
{-32'd1325, 32'd5970, -32'd917, -32'd280},
{-32'd15595, -32'd1714, 32'd1253, 32'd1246},
{-32'd5755, -32'd3724, 32'd5081, -32'd7020},
{-32'd22, -32'd5621, 32'd8427, 32'd9211},
{32'd348, 32'd3133, 32'd9422, -32'd325},
{-32'd9563, 32'd3866, 32'd7200, -32'd7758},
{32'd5693, -32'd3420, -32'd4348, 32'd4449},
{-32'd12628, 32'd5888, 32'd295, 32'd571},
{32'd5631, 32'd372, 32'd6434, -32'd10772},
{-32'd7720, 32'd5238, 32'd2177, 32'd3097},
{-32'd2954, 32'd2294, -32'd6346, -32'd2105},
{32'd2800, -32'd4485, 32'd1816, 32'd6289},
{32'd6450, 32'd5951, -32'd6497, 32'd6096},
{32'd3275, 32'd4097, -32'd2447, 32'd4144},
{32'd3727, -32'd8714, 32'd2694, 32'd847},
{-32'd1968, -32'd6160, 32'd4337, -32'd1055},
{-32'd6160, -32'd14365, -32'd3098, -32'd1904},
{32'd3595, -32'd2551, 32'd2241, -32'd582},
{32'd4904, 32'd1370, -32'd4039, 32'd9600},
{32'd4526, 32'd2160, 32'd894, 32'd8452},
{-32'd3789, -32'd1228, -32'd2137, 32'd9005},
{-32'd6189, -32'd7672, 32'd4884, -32'd7426},
{-32'd1198, 32'd6422, -32'd2304, 32'd1366},
{32'd1726, 32'd2826, 32'd8076, 32'd227},
{-32'd238, -32'd2321, 32'd3376, -32'd2961},
{-32'd7871, -32'd2548, -32'd4862, 32'd2705},
{-32'd2958, 32'd2476, -32'd2083, -32'd3763},
{-32'd12183, 32'd1593, 32'd5714, -32'd1276},
{-32'd6858, 32'd2936, 32'd3891, -32'd4963},
{32'd7700, -32'd5908, -32'd4652, -32'd3699},
{-32'd1351, -32'd6347, 32'd270, 32'd7016},
{-32'd2804, -32'd3160, -32'd2662, -32'd5798},
{32'd4841, 32'd5259, -32'd1658, 32'd5138},
{32'd3191, -32'd2537, -32'd4797, 32'd9552},
{-32'd8482, 32'd3526, 32'd3368, 32'd7817},
{-32'd4392, 32'd3322, 32'd2305, 32'd6685},
{-32'd10039, 32'd1268, -32'd2556, -32'd912},
{32'd5630, 32'd8176, -32'd6422, -32'd6422},
{-32'd4500, -32'd6212, 32'd3387, -32'd2538},
{-32'd3498, -32'd3524, -32'd5606, -32'd1426},
{-32'd459, -32'd9742, -32'd1525, 32'd4856},
{-32'd4, -32'd1453, -32'd1434, 32'd1635},
{-32'd4888, 32'd289, -32'd10153, -32'd3339},
{-32'd5932, -32'd1741, -32'd4344, -32'd2091},
{-32'd1977, 32'd2072, -32'd2208, 32'd4393},
{32'd439, 32'd1978, 32'd5244, -32'd855},
{32'd3184, -32'd93, 32'd6523, -32'd8243},
{-32'd11268, -32'd1580, -32'd2152, 32'd111},
{-32'd2478, 32'd1049, 32'd827, -32'd10005},
{32'd1236, 32'd7894, 32'd4819, 32'd3872},
{32'd3439, 32'd12430, 32'd8344, 32'd8744},
{-32'd3734, -32'd2055, -32'd3564, -32'd5216},
{32'd1389, -32'd5778, 32'd10188, -32'd203},
{32'd982, 32'd6659, -32'd7914, 32'd2363},
{-32'd10047, -32'd3744, -32'd63, -32'd3357},
{32'd6017, -32'd2138, 32'd8580, -32'd8812},
{32'd6257, -32'd4918, 32'd11361, -32'd994},
{32'd1648, -32'd5301, 32'd3755, -32'd4917},
{32'd1982, -32'd4622, 32'd5306, -32'd72},
{-32'd5787, -32'd5438, -32'd1498, -32'd4114},
{32'd3860, -32'd10037, -32'd3546, -32'd1337},
{-32'd5663, 32'd8282, -32'd8355, -32'd7002},
{-32'd1683, -32'd2803, -32'd5813, 32'd7198},
{32'd6305, 32'd8077, -32'd2909, 32'd1796},
{32'd540, -32'd3310, -32'd3109, 32'd2105},
{-32'd1853, 32'd11340, 32'd4208, 32'd8619},
{-32'd100, -32'd5878, 32'd3862, -32'd3753},
{32'd1954, 32'd483, 32'd5334, 32'd1267},
{-32'd11711, 32'd1774, -32'd2849, 32'd2693},
{-32'd1431, 32'd2675, 32'd5096, 32'd182},
{32'd193, -32'd7451, 32'd2733, -32'd11106},
{-32'd1033, 32'd586, -32'd8800, 32'd6642},
{32'd2919, -32'd1573, 32'd11310, 32'd4983},
{-32'd4492, -32'd49, -32'd4825, 32'd3119},
{-32'd1954, -32'd6498, -32'd9344, -32'd5836},
{-32'd278, -32'd6777, 32'd6483, -32'd2310},
{32'd6022, 32'd89, 32'd7141, -32'd8737},
{32'd5117, 32'd1012, -32'd7654, -32'd1725},
{32'd678, -32'd7100, 32'd9210, 32'd2319},
{32'd3143, -32'd3485, -32'd5530, 32'd1133},
{-32'd5641, 32'd5729, -32'd4896, -32'd6493},
{32'd1716, 32'd9209, -32'd2421, -32'd891},
{-32'd607, 32'd4740, -32'd10961, -32'd4976},
{32'd342, -32'd5689, 32'd2539, 32'd3844},
{-32'd1213, 32'd7205, -32'd1971, -32'd195},
{32'd6726, -32'd57, 32'd2223, 32'd2720},
{32'd4456, -32'd3117, 32'd2831, -32'd5378},
{-32'd4677, -32'd3282, -32'd3636, -32'd5932},
{-32'd2963, 32'd274, 32'd7186, 32'd1424},
{-32'd10428, 32'd1317, -32'd5607, -32'd1921},
{-32'd3242, -32'd4218, 32'd15087, -32'd3267},
{32'd7244, 32'd6205, -32'd1925, 32'd3584},
{32'd13004, -32'd917, -32'd5559, 32'd1338},
{-32'd194, 32'd4756, 32'd5271, 32'd4341},
{32'd1291, -32'd4638, -32'd10237, 32'd1869},
{32'd5352, -32'd440, -32'd6218, -32'd2436},
{32'd2860, -32'd1589, -32'd4928, -32'd1931},
{-32'd3138, -32'd1001, -32'd7346, -32'd4820},
{-32'd5314, -32'd5449, -32'd15527, 32'd1682},
{32'd6590, 32'd10621, 32'd7384, -32'd3193},
{32'd207, -32'd3268, -32'd8419, -32'd3826},
{-32'd3713, 32'd7055, 32'd787, -32'd2781},
{32'd2331, -32'd3385, 32'd5878, 32'd7970},
{32'd9919, 32'd5452, -32'd938, 32'd8022},
{-32'd7949, 32'd17762, -32'd3606, 32'd5730},
{-32'd7075, 32'd756, -32'd6902, 32'd1675},
{32'd8434, -32'd5583, 32'd8999, 32'd5710},
{32'd2610, 32'd2550, 32'd3467, 32'd489},
{32'd17646, -32'd7628, -32'd918, -32'd1353},
{-32'd6666, -32'd13126, 32'd1737, 32'd5973},
{32'd1940, -32'd6150, -32'd1347, 32'd2585},
{32'd8977, 32'd9355, 32'd3643, -32'd5198},
{32'd5273, -32'd4603, -32'd745, 32'd567},
{32'd9124, 32'd10140, 32'd1607, -32'd6499},
{-32'd9564, -32'd11191, 32'd5776, -32'd7759},
{32'd2764, -32'd13988, -32'd2102, -32'd1601},
{32'd5924, -32'd2060, -32'd5494, 32'd4108},
{32'd5615, -32'd7631, 32'd9772, 32'd5416},
{-32'd5726, -32'd12013, 32'd7182, -32'd1331},
{-32'd3017, 32'd4130, 32'd1412, -32'd8479},
{32'd2097, 32'd1265, -32'd4699, 32'd7106},
{32'd5874, 32'd1380, -32'd4719, 32'd268},
{-32'd5289, -32'd10249, -32'd9608, 32'd11689},
{32'd10733, 32'd2406, 32'd1736, 32'd2340},
{32'd3318, -32'd4450, 32'd7954, -32'd4906},
{-32'd4324, -32'd3696, 32'd7949, -32'd118},
{32'd1412, -32'd250, 32'd1408, 32'd562},
{-32'd7417, -32'd1405, -32'd7291, 32'd3607},
{32'd9737, 32'd5223, -32'd2031, 32'd4550},
{-32'd2358, 32'd11360, 32'd9448, 32'd8977},
{32'd2642, 32'd80, -32'd10851, 32'd6860},
{32'd1169, -32'd13096, 32'd9815, -32'd7121},
{-32'd2427, 32'd2146, -32'd3398, 32'd5163},
{32'd5374, 32'd8492, -32'd5325, -32'd217},
{-32'd2960, 32'd6583, 32'd7405, 32'd618},
{-32'd4471, 32'd4240, -32'd944, 32'd362},
{32'd80, -32'd11717, -32'd7766, -32'd1162},
{-32'd13618, 32'd4682, -32'd8094, 32'd6320},
{32'd9422, -32'd1839, 32'd588, 32'd56},
{32'd705, 32'd2925, -32'd3167, 32'd864},
{-32'd6508, -32'd6280, -32'd190, 32'd1874},
{32'd744, -32'd1863, 32'd3300, -32'd4399},
{32'd339, 32'd3423, -32'd453, -32'd4839},
{-32'd2852, -32'd2059, -32'd3755, -32'd3202},
{32'd103, 32'd5108, 32'd5049, 32'd1800},
{32'd3390, -32'd11, -32'd4330, -32'd2505},
{32'd3025, 32'd2046, -32'd10178, 32'd814}
},
{{32'd7429, -32'd6018, -32'd6792, -32'd1502},
{32'd8514, 32'd320, 32'd4264, 32'd8921},
{32'd1714, 32'd7224, 32'd5441, 32'd11804},
{32'd2621, 32'd4247, 32'd5629, -32'd7204},
{32'd7603, 32'd1355, 32'd8579, 32'd20025},
{-32'd8748, -32'd383, 32'd6485, 32'd465},
{32'd12231, -32'd873, 32'd5453, 32'd3831},
{32'd998, 32'd1354, -32'd9780, 32'd808},
{-32'd12987, 32'd6224, 32'd12005, -32'd5431},
{32'd9294, 32'd6994, 32'd7206, 32'd1822},
{-32'd2172, -32'd4802, 32'd98, 32'd5506},
{-32'd4290, 32'd1510, -32'd6189, 32'd3448},
{32'd6548, 32'd2257, 32'd6215, -32'd10716},
{32'd4513, 32'd5853, 32'd2051, 32'd1650},
{-32'd6175, -32'd14518, 32'd4655, -32'd8483},
{-32'd10220, -32'd11966, 32'd2010, -32'd5385},
{32'd6153, 32'd1759, 32'd2574, 32'd5316},
{-32'd4, 32'd3081, 32'd1993, 32'd2356},
{-32'd9151, -32'd8106, -32'd5537, 32'd4867},
{-32'd6334, 32'd1896, -32'd5093, 32'd5291},
{32'd738, 32'd10584, -32'd4883, -32'd6309},
{-32'd4601, -32'd2072, -32'd2377, -32'd1313},
{-32'd11702, -32'd1412, -32'd3905, -32'd1809},
{-32'd3876, -32'd4894, 32'd2564, -32'd3423},
{32'd4452, 32'd8128, 32'd1641, -32'd1208},
{32'd288, 32'd8263, 32'd12856, -32'd2880},
{-32'd10897, 32'd13280, -32'd2645, 32'd73},
{32'd1102, -32'd1052, 32'd2577, -32'd1723},
{32'd14878, 32'd16784, -32'd5070, 32'd1222},
{32'd4542, 32'd345, 32'd8092, 32'd1344},
{-32'd1593, -32'd7944, -32'd3456, 32'd8723},
{-32'd8990, -32'd10418, 32'd155, 32'd11881},
{32'd2858, 32'd1857, -32'd7402, 32'd5962},
{32'd1718, 32'd2769, 32'd3911, 32'd3241},
{32'd9717, 32'd1486, 32'd6760, -32'd1010},
{-32'd9328, -32'd13232, -32'd9968, 32'd5420},
{32'd5849, 32'd143, -32'd1753, -32'd3132},
{32'd3998, -32'd10840, 32'd9146, 32'd2836},
{32'd8446, 32'd206, -32'd6549, 32'd7405},
{32'd523, 32'd3924, 32'd4151, 32'd4416},
{32'd37, -32'd310, -32'd432, 32'd9580},
{32'd3038, -32'd5187, 32'd8428, 32'd2677},
{32'd7742, 32'd1762, 32'd9744, 32'd10812},
{-32'd1006, -32'd2879, 32'd4199, -32'd7960},
{-32'd1451, 32'd1729, -32'd10829, -32'd7415},
{32'd2615, -32'd8534, 32'd7901, -32'd4356},
{32'd4935, -32'd8263, -32'd1101, 32'd9756},
{-32'd3926, -32'd8784, -32'd6450, 32'd6779},
{-32'd2027, 32'd13318, -32'd2381, 32'd365},
{32'd2535, -32'd7716, -32'd3841, 32'd1214},
{-32'd430, 32'd8716, -32'd1767, 32'd7622},
{32'd7288, 32'd3407, 32'd1070, 32'd2523},
{32'd2524, 32'd5890, -32'd6663, 32'd4403},
{32'd1134, -32'd10338, 32'd17370, 32'd350},
{-32'd2733, -32'd196, 32'd5327, -32'd8661},
{-32'd2154, -32'd1690, -32'd11446, 32'd4191},
{-32'd4547, 32'd7989, -32'd7309, 32'd954},
{-32'd5947, -32'd12569, 32'd132, 32'd2315},
{-32'd4073, -32'd2471, -32'd1484, 32'd2359},
{-32'd3982, 32'd1876, -32'd1061, -32'd15542},
{32'd2282, -32'd3687, -32'd8193, -32'd6224},
{32'd1105, 32'd8480, -32'd11363, 32'd1583},
{-32'd5131, -32'd8278, 32'd119, 32'd5329},
{-32'd1465, -32'd3578, -32'd1689, -32'd5174},
{32'd1456, -32'd4803, 32'd1909, -32'd3586},
{32'd7812, 32'd9068, -32'd1687, 32'd3943},
{-32'd2651, -32'd6072, 32'd5847, -32'd6285},
{-32'd2488, 32'd4410, 32'd2154, -32'd4916},
{-32'd1795, -32'd4515, -32'd15977, -32'd5191},
{-32'd3911, -32'd6649, -32'd1620, -32'd667},
{32'd1409, -32'd11040, -32'd1405, 32'd2248},
{32'd12170, 32'd6280, 32'd11385, 32'd5678},
{-32'd4770, -32'd3649, -32'd4371, -32'd2886},
{32'd527, -32'd1538, -32'd8135, -32'd4028},
{32'd228, 32'd4878, -32'd2718, -32'd9865},
{32'd893, -32'd413, 32'd1992, -32'd4442},
{32'd1101, 32'd4990, 32'd844, 32'd7783},
{-32'd5817, -32'd3227, -32'd383, 32'd633},
{32'd8451, 32'd7689, 32'd4621, -32'd1471},
{32'd3485, 32'd8565, 32'd2745, 32'd2588},
{32'd6415, -32'd2841, -32'd5751, -32'd6528},
{32'd1419, -32'd2686, -32'd5452, 32'd8269},
{-32'd2470, 32'd3977, -32'd10164, 32'd630},
{32'd6877, -32'd120, 32'd3294, 32'd9289},
{-32'd4271, 32'd1377, -32'd9328, 32'd7549},
{32'd1871, -32'd4906, 32'd8059, 32'd6591},
{32'd599, -32'd7334, 32'd8625, 32'd3876},
{-32'd4579, -32'd10533, -32'd4247, -32'd4140},
{32'd2074, 32'd4261, 32'd9704, 32'd422},
{32'd3668, -32'd9853, -32'd994, 32'd7452},
{32'd14211, 32'd1591, 32'd4266, -32'd6813},
{-32'd3113, -32'd10701, -32'd5691, 32'd6542},
{32'd5624, -32'd514, 32'd8277, 32'd3026},
{32'd3878, 32'd6762, 32'd8416, 32'd4504},
{32'd18291, 32'd6996, -32'd1585, 32'd5051},
{32'd1311, 32'd7308, 32'd37, 32'd7977},
{32'd1866, 32'd683, -32'd9707, 32'd7219},
{-32'd1305, 32'd782, 32'd5898, -32'd5298},
{32'd9183, 32'd826, 32'd6669, 32'd1203},
{32'd3782, 32'd1532, 32'd6300, 32'd1631},
{-32'd1192, -32'd16178, -32'd4556, -32'd5593},
{32'd1811, -32'd3347, -32'd4502, 32'd6407},
{-32'd831, 32'd10900, 32'd6859, 32'd4776},
{-32'd3010, 32'd11035, -32'd7551, 32'd2432},
{32'd8297, -32'd6608, -32'd9194, 32'd904},
{-32'd1515, -32'd5640, -32'd1505, 32'd805},
{-32'd1702, 32'd2780, 32'd2541, 32'd63},
{-32'd10057, -32'd4394, -32'd16304, 32'd3145},
{-32'd6612, -32'd5169, -32'd1162, -32'd13912},
{-32'd6661, -32'd4539, -32'd213, -32'd5827},
{-32'd424, 32'd442, -32'd12672, -32'd4616},
{32'd1829, 32'd2558, -32'd2309, 32'd3520},
{32'd1147, -32'd2980, 32'd9000, 32'd5833},
{-32'd3452, -32'd4083, -32'd685, 32'd5339},
{-32'd8035, -32'd10207, 32'd2850, -32'd4060},
{-32'd637, -32'd8387, -32'd7107, -32'd13691},
{-32'd2237, 32'd39, -32'd4901, 32'd527},
{-32'd6107, 32'd7439, -32'd4528, -32'd3889},
{32'd3712, 32'd4795, 32'd7976, 32'd713},
{-32'd5823, -32'd2364, 32'd4897, 32'd1666},
{-32'd5782, 32'd2866, 32'd3243, 32'd1702},
{32'd834, -32'd695, -32'd3626, -32'd4310},
{32'd102, 32'd2089, 32'd2142, 32'd989},
{-32'd1199, 32'd9220, 32'd5860, 32'd1626},
{-32'd829, -32'd9329, -32'd9389, 32'd6513},
{32'd5051, 32'd9741, 32'd8275, -32'd11428},
{-32'd6869, -32'd5090, -32'd8150, -32'd5812},
{-32'd12728, 32'd1543, -32'd1876, -32'd4951},
{32'd1121, -32'd10364, 32'd121, -32'd3292},
{-32'd5377, 32'd2582, -32'd6303, 32'd2835},
{-32'd4321, -32'd10038, -32'd15646, -32'd2668},
{32'd14590, -32'd2794, -32'd435, 32'd9914},
{-32'd10534, -32'd1778, -32'd16179, -32'd9340},
{32'd6266, 32'd11674, 32'd3997, 32'd8398},
{-32'd3796, 32'd779, 32'd4808, -32'd5756},
{32'd10940, -32'd7803, -32'd8110, 32'd5454},
{32'd7335, -32'd107, 32'd3483, 32'd2053},
{-32'd6635, -32'd3019, 32'd4394, -32'd476},
{32'd13730, 32'd14257, 32'd8007, -32'd3940},
{32'd5000, -32'd3484, -32'd14428, -32'd5857},
{-32'd799, -32'd6843, -32'd7718, 32'd650},
{32'd7918, 32'd8373, -32'd761, 32'd13313},
{-32'd6424, -32'd3423, -32'd3293, 32'd3492},
{32'd11268, 32'd1661, -32'd4955, 32'd220},
{32'd2148, 32'd6830, -32'd5120, 32'd546},
{32'd6526, 32'd2256, 32'd12084, -32'd3045},
{-32'd664, -32'd507, -32'd704, -32'd716},
{32'd1025, -32'd10106, 32'd8382, -32'd4185},
{-32'd3256, 32'd8654, 32'd7210, 32'd825},
{-32'd7096, 32'd2592, 32'd238, 32'd997},
{32'd1289, -32'd2020, 32'd4783, 32'd4192},
{32'd1634, 32'd3486, 32'd2141, 32'd2116},
{-32'd3118, 32'd10262, -32'd4825, -32'd8656},
{32'd5172, 32'd4076, 32'd6419, 32'd761},
{32'd1393, -32'd10027, 32'd285, 32'd4222},
{32'd6803, -32'd5231, 32'd6075, -32'd6051},
{-32'd4160, 32'd2706, 32'd4791, -32'd3082},
{32'd7127, -32'd60, -32'd137, -32'd4372},
{-32'd2748, -32'd2098, 32'd4480, -32'd4064},
{32'd5396, 32'd8080, -32'd8516, 32'd478},
{-32'd13385, -32'd8484, -32'd9162, -32'd7143},
{32'd2167, 32'd15332, -32'd2203, -32'd1998},
{-32'd9184, 32'd2350, -32'd10701, 32'd843},
{32'd12589, 32'd10469, 32'd9583, 32'd3305},
{32'd5412, 32'd12915, 32'd11359, 32'd2868},
{-32'd4807, -32'd10131, 32'd3336, 32'd2917},
{32'd966, 32'd2712, 32'd9265, 32'd8300},
{-32'd3014, -32'd3266, -32'd13542, -32'd458},
{32'd10577, -32'd12467, -32'd21, 32'd6553},
{-32'd15193, -32'd11170, -32'd10390, 32'd3582},
{-32'd5421, -32'd16736, 32'd7105, 32'd11707},
{-32'd1227, -32'd2580, -32'd3335, -32'd10174},
{32'd9275, -32'd565, 32'd6523, -32'd5959},
{-32'd10981, -32'd1000, -32'd416, 32'd2717},
{-32'd4778, 32'd13517, 32'd13284, 32'd4735},
{32'd3341, -32'd15603, -32'd6476, 32'd14727},
{-32'd3729, 32'd9364, -32'd6609, 32'd754},
{32'd5539, 32'd6726, 32'd2651, 32'd2429},
{-32'd4569, -32'd8897, -32'd4724, 32'd2885},
{-32'd2039, -32'd7586, 32'd86, 32'd4046},
{-32'd7358, -32'd1181, -32'd5839, 32'd3982},
{-32'd1037, -32'd4049, -32'd4044, -32'd5793},
{-32'd7757, 32'd8667, -32'd1538, 32'd3081},
{32'd12080, -32'd13897, 32'd4234, -32'd5649},
{32'd984, 32'd147, 32'd4447, -32'd387},
{-32'd3438, -32'd451, -32'd10100, 32'd768},
{-32'd4378, 32'd10948, 32'd5058, 32'd1470},
{32'd5490, -32'd9714, -32'd386, -32'd4905},
{32'd3629, 32'd1667, 32'd12176, -32'd12291},
{32'd604, -32'd7571, -32'd2017, -32'd7108},
{32'd5737, -32'd2099, 32'd4618, 32'd2069},
{-32'd5302, -32'd1005, 32'd5280, -32'd4018},
{-32'd15, 32'd3979, 32'd8688, -32'd11432},
{32'd3736, 32'd791, 32'd7658, -32'd4656},
{32'd4568, -32'd2139, 32'd755, -32'd2071},
{-32'd9326, -32'd2427, -32'd16767, -32'd2171},
{-32'd4624, -32'd7369, -32'd1222, 32'd6310},
{32'd90, 32'd5319, -32'd8912, 32'd4584},
{32'd4588, -32'd10548, -32'd10378, 32'd5812},
{-32'd2982, -32'd17, -32'd2831, 32'd2302},
{-32'd5381, -32'd9561, -32'd9926, 32'd904},
{32'd10713, -32'd1441, 32'd5453, 32'd471},
{-32'd4939, 32'd1763, -32'd4772, 32'd6339},
{32'd7131, 32'd9227, 32'd9463, 32'd1244},
{32'd2211, -32'd2581, -32'd7017, 32'd6546},
{-32'd3233, -32'd2441, 32'd8748, -32'd3066},
{32'd1679, -32'd4426, -32'd14887, -32'd3346},
{-32'd4036, -32'd204, 32'd4285, -32'd6982},
{32'd6166, 32'd611, 32'd3663, -32'd5166},
{32'd6625, 32'd11806, 32'd3736, 32'd2255},
{32'd15999, -32'd5603, 32'd4818, -32'd3180},
{-32'd466, -32'd1949, -32'd3576, 32'd710},
{32'd6353, -32'd5991, 32'd8497, -32'd3745},
{-32'd8758, 32'd766, 32'd9262, 32'd8119},
{32'd2620, 32'd2239, 32'd1266, -32'd3775},
{-32'd3835, -32'd5976, 32'd2642, 32'd3664},
{32'd678, -32'd8185, 32'd7097, -32'd9672},
{-32'd1934, -32'd3031, 32'd10499, -32'd4479},
{-32'd385, 32'd3420, 32'd6492, -32'd916},
{32'd3522, 32'd3784, 32'd2249, 32'd510},
{32'd5031, -32'd3694, 32'd10807, 32'd6088},
{32'd1101, 32'd11613, 32'd1591, -32'd7459},
{32'd12498, 32'd17534, -32'd6617, -32'd10653},
{-32'd6196, 32'd7311, -32'd1200, 32'd8395},
{-32'd1165, 32'd4660, -32'd254, 32'd372},
{32'd3902, 32'd3230, 32'd2179, -32'd769},
{32'd2785, -32'd8425, 32'd4638, -32'd2572},
{-32'd5637, 32'd4609, -32'd8138, -32'd2393},
{32'd2233, 32'd4041, -32'd9682, -32'd958},
{32'd3492, 32'd627, -32'd180, -32'd7587},
{-32'd4370, -32'd12499, -32'd5198, 32'd2642},
{-32'd820, 32'd9124, 32'd138, -32'd1861},
{32'd5626, -32'd11106, 32'd3853, -32'd1403},
{32'd6364, 32'd8278, -32'd2614, 32'd3430},
{-32'd6778, -32'd2325, 32'd8371, 32'd8269},
{32'd178, -32'd1554, 32'd3509, -32'd7339},
{-32'd9725, -32'd6591, -32'd1314, 32'd9733},
{32'd2278, -32'd4151, 32'd5782, 32'd3932},
{32'd871, 32'd5159, 32'd6472, 32'd2554},
{-32'd103, -32'd2777, 32'd2953, 32'd2091},
{-32'd7306, -32'd4453, -32'd8659, 32'd3011},
{32'd10901, -32'd6113, 32'd2473, 32'd6977},
{-32'd9380, 32'd2941, -32'd864, 32'd3084},
{-32'd24, -32'd3005, 32'd7717, -32'd5236},
{32'd9512, 32'd552, -32'd621, -32'd4232},
{-32'd6539, -32'd1566, -32'd10507, -32'd10675},
{32'd3471, -32'd16781, 32'd352, 32'd6537},
{-32'd3067, -32'd2042, 32'd505, 32'd11384},
{32'd2188, -32'd4797, 32'd4623, 32'd4712},
{-32'd412, 32'd2252, 32'd6183, -32'd2646},
{32'd8024, -32'd11492, 32'd4962, -32'd6222},
{-32'd5549, 32'd30, -32'd4906, 32'd9397},
{32'd6031, 32'd14001, 32'd5076, -32'd6507},
{-32'd10366, -32'd5232, -32'd1763, -32'd1416},
{32'd1694, -32'd579, -32'd7400, 32'd535},
{-32'd7215, -32'd3264, 32'd12429, 32'd10482},
{32'd768, 32'd8514, -32'd11475, 32'd5609},
{32'd10227, 32'd9578, 32'd1101, -32'd10340},
{-32'd4135, -32'd13213, -32'd9222, -32'd776},
{-32'd6637, 32'd5133, 32'd6592, -32'd3901},
{-32'd1169, -32'd2168, -32'd555, -32'd11638},
{32'd1648, 32'd3826, 32'd10983, -32'd6286},
{-32'd2492, 32'd159, -32'd1752, 32'd5369},
{32'd16433, -32'd4380, -32'd8274, -32'd393},
{32'd1801, 32'd12864, 32'd1837, 32'd1872},
{-32'd920, -32'd3275, -32'd8082, 32'd2709},
{-32'd5026, -32'd1488, -32'd3288, -32'd3467},
{-32'd4946, -32'd6477, -32'd3834, 32'd14355},
{-32'd426, -32'd2485, 32'd2359, 32'd821},
{-32'd8604, -32'd6696, -32'd1135, 32'd12948},
{-32'd591, -32'd6185, 32'd4498, -32'd9200},
{-32'd285, -32'd6436, 32'd7734, -32'd13106},
{32'd5300, -32'd1250, -32'd3873, 32'd11318},
{-32'd2648, -32'd385, 32'd9108, 32'd6521},
{32'd3201, -32'd5869, -32'd5793, 32'd4218},
{-32'd4532, 32'd2514, 32'd4817, 32'd8444},
{32'd10957, 32'd4231, 32'd5297, 32'd300},
{-32'd15885, 32'd10716, 32'd5773, 32'd5350},
{-32'd12573, -32'd2252, -32'd3782, -32'd5757},
{32'd1320, -32'd10658, -32'd3389, 32'd3887},
{32'd7910, -32'd565, -32'd656, -32'd3894},
{32'd11608, -32'd8004, 32'd2433, -32'd5586},
{32'd7465, -32'd5717, 32'd862, -32'd574},
{-32'd4479, -32'd2207, 32'd5093, 32'd2456},
{-32'd6720, 32'd1865, -32'd8157, 32'd831},
{-32'd5746, -32'd10510, -32'd5328, 32'd7750},
{-32'd4508, 32'd1833, -32'd166, -32'd7570},
{-32'd9619, -32'd9568, 32'd683, -32'd5190},
{32'd1926, 32'd2153, 32'd6426, 32'd14906},
{-32'd2516, -32'd14540, -32'd2103, 32'd1250},
{32'd2180, 32'd399, -32'd2745, -32'd8251},
{32'd7678, 32'd15769, -32'd871, -32'd6834},
{-32'd849, -32'd204, -32'd9553, -32'd1054},
{32'd5818, -32'd12799, -32'd15386, 32'd12246},
{32'd2506, -32'd8175, -32'd5763, -32'd2593},
{-32'd979, -32'd4962, 32'd7953, 32'd4682},
{-32'd102, 32'd10, -32'd3680, -32'd6400},
{-32'd1362, 32'd960, -32'd2626, 32'd1216},
{-32'd6314, 32'd1919, 32'd564, -32'd9224},
{-32'd10820, -32'd10904, -32'd8881, 32'd4349}
},
{{32'd12641, 32'd12669, 32'd9003, 32'd326},
{-32'd4463, -32'd991, 32'd9300, -32'd7777},
{-32'd2382, 32'd2392, 32'd8878, -32'd9604},
{32'd5589, 32'd7110, 32'd2317, 32'd2352},
{-32'd11064, 32'd2947, -32'd2934, 32'd4454},
{32'd730, -32'd5488, 32'd3458, -32'd2831},
{32'd14224, -32'd4190, 32'd2912, -32'd872},
{32'd991, -32'd7387, 32'd7060, -32'd5180},
{-32'd6241, 32'd3533, -32'd7066, -32'd7322},
{32'd12622, 32'd1720, 32'd5366, 32'd6129},
{-32'd2219, 32'd4107, 32'd1419, -32'd8451},
{32'd4608, 32'd7794, -32'd4865, 32'd3641},
{32'd3437, -32'd2902, 32'd9780, 32'd3940},
{-32'd8763, -32'd16875, -32'd2305, -32'd4043},
{-32'd3659, -32'd3317, -32'd16024, -32'd118},
{32'd1573, -32'd807, -32'd2691, -32'd2375},
{32'd2473, -32'd14, 32'd3584, 32'd5157},
{32'd1577, 32'd2921, 32'd9780, -32'd5375},
{32'd3355, -32'd3847, -32'd6957, -32'd1872},
{32'd6293, -32'd2906, 32'd1528, 32'd4382},
{32'd4431, 32'd2033, -32'd928, 32'd3973},
{-32'd8342, -32'd4855, -32'd1064, 32'd1699},
{-32'd8116, -32'd14, -32'd4531, -32'd431},
{-32'd1573, -32'd7866, -32'd2621, 32'd3140},
{32'd7449, -32'd4708, 32'd12818, -32'd2166},
{-32'd3507, 32'd8308, -32'd2735, -32'd6642},
{-32'd4134, -32'd279, -32'd3590, -32'd4902},
{-32'd3628, -32'd2078, -32'd270, -32'd5196},
{32'd4515, 32'd478, 32'd12527, -32'd87},
{-32'd4916, -32'd2440, -32'd3830, -32'd3106},
{-32'd6284, -32'd2911, -32'd3996, 32'd110},
{-32'd10889, -32'd6500, 32'd650, -32'd3939},
{32'd14422, 32'd9313, 32'd4951, 32'd3630},
{-32'd13889, 32'd2306, -32'd4486, -32'd612},
{32'd10300, -32'd1644, 32'd6027, 32'd6034},
{-32'd2765, 32'd3997, 32'd5275, -32'd2489},
{32'd1548, 32'd5477, -32'd2329, 32'd4891},
{32'd4868, 32'd10313, -32'd3641, 32'd3929},
{32'd11681, 32'd9222, -32'd5906, -32'd2957},
{32'd7666, -32'd1262, -32'd12489, 32'd7741},
{32'd11989, -32'd3171, 32'd446, -32'd1639},
{32'd1872, 32'd7085, 32'd5661, -32'd1401},
{-32'd3691, -32'd5362, 32'd1086, 32'd4032},
{-32'd8501, -32'd14529, -32'd8008, 32'd1193},
{-32'd5394, 32'd1933, -32'd10970, -32'd821},
{-32'd5312, -32'd3886, 32'd3484, -32'd5097},
{32'd3088, -32'd13329, -32'd590, -32'd1365},
{-32'd6114, -32'd8266, -32'd3363, 32'd3174},
{32'd9887, 32'd10832, 32'd5459, 32'd1361},
{32'd5863, 32'd6124, 32'd5336, -32'd7459},
{32'd6060, -32'd5038, -32'd138, -32'd2476},
{32'd3489, 32'd3957, 32'd4405, -32'd1948},
{-32'd3759, 32'd2154, 32'd4040, -32'd580},
{32'd8180, 32'd7606, -32'd6814, -32'd5389},
{32'd10449, 32'd6202, 32'd6013, 32'd8991},
{-32'd10192, 32'd1198, -32'd3509, -32'd7574},
{32'd7593, -32'd1579, -32'd448, -32'd11},
{-32'd13578, -32'd4499, -32'd2617, -32'd9070},
{-32'd3947, -32'd2095, -32'd9933, -32'd5969},
{32'd4849, 32'd3635, 32'd2980, -32'd3967},
{-32'd9246, -32'd956, -32'd1509, -32'd2684},
{32'd9519, 32'd2572, -32'd4502, 32'd1606},
{-32'd5667, -32'd2473, -32'd2145, -32'd4611},
{-32'd12532, -32'd667, -32'd6664, 32'd694},
{32'd185, 32'd5544, -32'd531, -32'd1439},
{32'd6377, 32'd3608, 32'd12633, 32'd593},
{32'd1546, -32'd4206, -32'd11678, 32'd1114},
{-32'd559, -32'd1629, -32'd2977, -32'd5308},
{-32'd1549, -32'd5178, 32'd13481, 32'd1496},
{-32'd188, -32'd1741, -32'd1112, -32'd1903},
{-32'd5591, 32'd73, -32'd10615, -32'd5195},
{-32'd8818, 32'd20, 32'd1842, -32'd3388},
{-32'd12469, 32'd897, -32'd989, 32'd265},
{32'd7743, -32'd996, -32'd4067, 32'd4348},
{32'd2485, 32'd6265, 32'd548, -32'd2063},
{32'd1401, -32'd2823, 32'd259, -32'd2479},
{-32'd8335, -32'd7946, -32'd2316, -32'd4646},
{-32'd493, 32'd5665, -32'd7628, -32'd5353},
{32'd12718, 32'd5841, 32'd15246, 32'd4422},
{32'd641, 32'd2022, -32'd7646, -32'd1114},
{32'd11701, 32'd239, 32'd78, 32'd4590},
{32'd36, -32'd1362, 32'd13429, -32'd782},
{-32'd12562, -32'd2997, -32'd2473, -32'd5906},
{-32'd2222, 32'd6863, -32'd344, 32'd1670},
{-32'd10138, -32'd1622, 32'd8318, -32'd6561},
{-32'd4483, -32'd3103, -32'd6428, -32'd3480},
{32'd9821, 32'd10166, 32'd6358, 32'd7152},
{-32'd4884, -32'd2220, -32'd10105, -32'd2411},
{-32'd1688, -32'd3755, 32'd2144, -32'd11200},
{-32'd8776, -32'd3022, -32'd75, -32'd1983},
{32'd10829, 32'd67, 32'd12779, 32'd2673},
{-32'd8365, -32'd1094, -32'd8900, -32'd1221},
{-32'd2323, 32'd1187, -32'd9170, 32'd7933},
{32'd1368, 32'd2729, 32'd3628, -32'd2123},
{-32'd3845, 32'd4111, 32'd914, -32'd4306},
{-32'd5225, -32'd1996, 32'd3643, -32'd3096},
{32'd4869, 32'd918, 32'd1150, 32'd5673},
{-32'd11247, 32'd1911, 32'd4067, -32'd1326},
{-32'd3007, 32'd1850, -32'd1837, -32'd2058},
{32'd9463, 32'd5867, 32'd3588, 32'd10169},
{-32'd7036, -32'd4229, -32'd3246, -32'd620},
{-32'd10713, -32'd1913, 32'd5403, -32'd8634},
{-32'd1296, -32'd1461, 32'd5483, 32'd4907},
{32'd5928, 32'd10094, 32'd8259, 32'd2307},
{-32'd2831, 32'd383, 32'd7961, 32'd8399},
{-32'd3391, -32'd3669, -32'd11340, -32'd4665},
{-32'd8983, -32'd9158, -32'd2187, -32'd5451},
{-32'd4202, 32'd167, -32'd8870, 32'd1045},
{32'd2185, 32'd1898, 32'd1862, 32'd7686},
{-32'd12628, -32'd5953, -32'd12980, -32'd573},
{-32'd1206, 32'd1818, -32'd4440, 32'd926},
{32'd2551, 32'd2028, 32'd4203, 32'd2265},
{32'd10385, 32'd4119, 32'd6619, 32'd4515},
{32'd3487, 32'd8192, 32'd13328, 32'd2853},
{-32'd3998, -32'd463, -32'd5763, -32'd3190},
{32'd827, -32'd1146, 32'd2642, -32'd2379},
{32'd4581, 32'd64, 32'd2741, 32'd4025},
{-32'd7769, -32'd6410, 32'd11618, 32'd2036},
{-32'd569, 32'd1240, 32'd1492, -32'd1731},
{32'd8908, 32'd4470, -32'd2592, 32'd1176},
{32'd13484, 32'd3216, -32'd3219, 32'd3198},
{32'd1890, 32'd7067, -32'd12154, -32'd1307},
{32'd3497, -32'd5925, 32'd2883, -32'd2634},
{-32'd3689, -32'd8563, -32'd3379, -32'd3430},
{-32'd6258, -32'd2135, 32'd3268, 32'd2535},
{-32'd1624, -32'd4362, 32'd3531, 32'd4529},
{32'd4007, 32'd7992, -32'd10395, 32'd649},
{-32'd6781, -32'd9541, -32'd5903, -32'd4233},
{-32'd2681, 32'd3343, -32'd11898, 32'd2005},
{32'd9230, 32'd3050, -32'd1083, -32'd2563},
{-32'd1734, -32'd3777, -32'd3233, 32'd2997},
{32'd1604, 32'd1298, 32'd9047, -32'd2693},
{-32'd2692, -32'd7483, -32'd13216, 32'd3442},
{-32'd4219, -32'd3197, 32'd8478, -32'd6300},
{-32'd7823, -32'd14997, 32'd146, -32'd320},
{-32'd17777, -32'd3412, -32'd6104, -32'd5885},
{-32'd16153, -32'd9280, 32'd5852, -32'd2522},
{32'd8659, 32'd3184, -32'd6269, -32'd6064},
{32'd838, 32'd3837, 32'd4528, -32'd93},
{32'd6220, -32'd2019, 32'd4760, -32'd5141},
{32'd7264, 32'd2645, -32'd3950, 32'd3106},
{-32'd4487, -32'd5287, 32'd3645, -32'd518},
{-32'd2493, 32'd8387, -32'd3449, -32'd2014},
{-32'd6530, -32'd3777, 32'd11348, -32'd3394},
{32'd2173, 32'd4557, 32'd2845, 32'd8458},
{32'd1657, 32'd11236, 32'd11655, -32'd5206},
{-32'd7805, -32'd2712, -32'd6919, 32'd1844},
{32'd15, -32'd7293, -32'd8674, 32'd5054},
{32'd5256, -32'd4807, 32'd4623, -32'd2911},
{-32'd2688, -32'd16485, -32'd5931, -32'd1064},
{32'd2125, 32'd6181, -32'd782, 32'd335},
{-32'd6147, 32'd6850, 32'd9089, 32'd2726},
{-32'd4025, 32'd6730, 32'd3603, 32'd1832},
{32'd1702, -32'd3374, 32'd2130, 32'd7373},
{-32'd9400, -32'd11115, 32'd1602, 32'd1780},
{-32'd5917, 32'd3526, -32'd19586, 32'd531},
{32'd1472, 32'd2566, 32'd1465, 32'd2661},
{32'd6987, 32'd1242, 32'd2035, -32'd8442},
{-32'd5236, 32'd6514, -32'd13574, 32'd5609},
{-32'd1802, -32'd3332, -32'd1897, 32'd1955},
{-32'd12775, 32'd576, 32'd301, -32'd14229},
{32'd6712, 32'd4650, 32'd2863, 32'd1327},
{-32'd11810, -32'd4547, -32'd5113, 32'd2807},
{32'd7286, 32'd8525, 32'd9471, 32'd4648},
{-32'd2663, 32'd1746, 32'd10213, 32'd3697},
{32'd2245, -32'd3581, -32'd2974, -32'd2593},
{-32'd8253, -32'd10258, -32'd825, 32'd2211},
{-32'd2701, -32'd566, -32'd6388, -32'd7484},
{32'd4149, 32'd981, 32'd2689, -32'd1967},
{32'd2479, -32'd68, -32'd7715, -32'd1558},
{-32'd5180, -32'd970, -32'd3847, 32'd990},
{-32'd6354, -32'd6863, -32'd9564, 32'd659},
{32'd2814, -32'd1300, 32'd7850, 32'd4602},
{32'd2489, 32'd6260, -32'd941, 32'd840},
{-32'd7043, 32'd1352, -32'd168, 32'd9448},
{32'd2049, 32'd1848, -32'd1872, 32'd5707},
{32'd2689, 32'd723, -32'd4341, 32'd617},
{32'd1243, 32'd6192, 32'd204, -32'd8370},
{-32'd5205, -32'd6822, 32'd2999, 32'd856},
{32'd94, -32'd3164, -32'd2728, -32'd2329},
{-32'd7690, 32'd277, 32'd3369, 32'd4181},
{32'd7764, 32'd358, -32'd2617, -32'd434},
{32'd2577, 32'd3541, 32'd1529, -32'd7960},
{-32'd3386, -32'd1017, 32'd6024, 32'd50},
{-32'd1614, -32'd2835, 32'd5585, 32'd6565},
{32'd7745, 32'd5330, -32'd2622, 32'd392},
{32'd531, -32'd4613, 32'd10897, -32'd2972},
{32'd2072, 32'd4249, -32'd5645, 32'd3379},
{-32'd9075, -32'd6495, -32'd163, 32'd932},
{-32'd6284, -32'd3542, 32'd5521, -32'd1822},
{32'd3322, 32'd3731, -32'd3995, 32'd4132},
{-32'd6649, -32'd6031, -32'd3696, -32'd2573},
{-32'd9812, 32'd7197, -32'd9242, -32'd4785},
{-32'd6204, -32'd11751, 32'd4532, 32'd6907},
{32'd6312, -32'd7830, -32'd1256, -32'd9931},
{-32'd1627, -32'd102, -32'd347, 32'd2495},
{-32'd11029, -32'd2294, -32'd2145, 32'd4465},
{32'd2574, 32'd8459, 32'd2026, -32'd2060},
{32'd8699, 32'd3874, 32'd10604, 32'd548},
{32'd3553, 32'd9229, 32'd93, -32'd4452},
{-32'd3522, -32'd6010, -32'd3335, -32'd2765},
{-32'd3378, 32'd129, -32'd8844, -32'd1995},
{32'd4983, 32'd7378, 32'd8017, 32'd6881},
{32'd3159, 32'd4085, 32'd8262, 32'd451},
{-32'd10268, 32'd3074, 32'd4031, -32'd578},
{-32'd10599, -32'd5183, 32'd1532, 32'd5052},
{32'd8666, 32'd3584, -32'd2347, -32'd333},
{-32'd3526, -32'd54, 32'd57, 32'd2299},
{32'd1966, -32'd8705, 32'd5863, -32'd949},
{32'd2486, -32'd2594, 32'd7010, -32'd4645},
{32'd797, 32'd4652, 32'd1992, -32'd623},
{32'd2203, 32'd298, -32'd3820, -32'd2528},
{32'd380, 32'd11876, 32'd1241, 32'd3136},
{-32'd5146, 32'd7660, -32'd9846, -32'd5783},
{32'd1171, 32'd9266, 32'd2617, 32'd168},
{32'd2512, -32'd9964, -32'd3426, 32'd3180},
{-32'd1741, -32'd12362, 32'd10584, -32'd1102},
{-32'd4602, -32'd25, 32'd3487, 32'd4203},
{-32'd3030, 32'd3036, 32'd6278, 32'd10449},
{-32'd6789, 32'd200, 32'd6228, -32'd1521},
{-32'd9771, -32'd10052, 32'd6483, -32'd4685},
{32'd4616, 32'd5094, 32'd2310, 32'd638},
{32'd11744, -32'd4692, -32'd7397, 32'd834},
{-32'd3553, -32'd13448, -32'd2921, -32'd4385},
{-32'd4499, -32'd1909, 32'd1283, 32'd5632},
{32'd3473, -32'd8960, 32'd10798, 32'd4276},
{-32'd3190, -32'd4536, 32'd10552, 32'd1814},
{32'd2571, 32'd2001, -32'd3607, -32'd7854},
{32'd12575, -32'd10266, 32'd10507, -32'd4540},
{32'd2713, 32'd5635, -32'd1200, 32'd1100},
{-32'd138, -32'd7520, -32'd5312, -32'd3891},
{-32'd12291, -32'd1469, -32'd12244, 32'd242},
{32'd694, 32'd1694, 32'd2474, -32'd2130},
{-32'd3452, 32'd5518, -32'd4183, -32'd1151},
{-32'd5832, -32'd6743, -32'd35, -32'd1079},
{-32'd10555, -32'd6328, 32'd5516, -32'd746},
{32'd5403, 32'd596, 32'd5060, -32'd943},
{-32'd8447, 32'd5587, 32'd5829, -32'd1926},
{32'd1227, 32'd5898, -32'd7172, 32'd3887},
{-32'd1228, -32'd2018, -32'd1787, 32'd109},
{-32'd779, 32'd9920, -32'd4526, 32'd3527},
{-32'd9535, -32'd498, -32'd5436, -32'd7398},
{-32'd7658, -32'd9610, -32'd9320, 32'd614},
{32'd1486, -32'd1232, -32'd230, 32'd2068},
{32'd6039, 32'd6981, -32'd815, 32'd5294},
{-32'd2910, 32'd160, -32'd15182, 32'd1795},
{-32'd1556, -32'd6915, 32'd2232, 32'd3097},
{32'd682, -32'd10499, -32'd2373, -32'd1466},
{32'd126, -32'd1708, 32'd4594, 32'd2014},
{32'd997, 32'd2058, -32'd4637, -32'd2133},
{-32'd1488, 32'd3327, 32'd3109, -32'd627},
{-32'd4445, -32'd11110, 32'd1165, -32'd1949},
{-32'd2126, 32'd8275, 32'd6718, -32'd2300},
{32'd11093, -32'd7659, 32'd5234, 32'd6959},
{-32'd5791, -32'd1288, 32'd4834, -32'd1977},
{-32'd6443, -32'd5142, -32'd585, 32'd2279},
{32'd8356, -32'd257, -32'd6944, 32'd4399},
{32'd8396, 32'd3563, 32'd6529, 32'd13422},
{32'd2490, 32'd6187, -32'd2124, -32'd1405},
{32'd6611, 32'd2375, -32'd304, 32'd8512},
{-32'd1745, -32'd8608, -32'd2400, 32'd4623},
{-32'd2323, 32'd986, -32'd12825, -32'd6457},
{32'd4461, 32'd4596, 32'd2470, 32'd1995},
{-32'd1216, 32'd3281, -32'd7291, 32'd7967},
{32'd3487, 32'd5051, -32'd4086, 32'd1696},
{-32'd5846, -32'd2742, -32'd3732, -32'd7325},
{32'd10749, 32'd8026, -32'd6359, 32'd5229},
{-32'd2273, 32'd9823, -32'd7564, -32'd3087},
{-32'd321, -32'd2026, 32'd5703, -32'd1969},
{-32'd7323, 32'd3255, 32'd763, -32'd9155},
{-32'd10, -32'd3080, 32'd2829, -32'd4453},
{32'd4126, 32'd4265, -32'd390, -32'd4154},
{-32'd6229, -32'd10101, 32'd5911, 32'd1785},
{-32'd7046, -32'd14293, 32'd3544, -32'd401},
{32'd9345, 32'd1336, -32'd1090, -32'd6086},
{32'd6626, -32'd1763, -32'd3899, -32'd6616},
{32'd11803, 32'd6112, 32'd4925, 32'd5412},
{-32'd9190, 32'd3274, 32'd709, -32'd1563},
{-32'd6159, 32'd3222, -32'd14019, -32'd2022},
{32'd2860, -32'd297, -32'd13955, -32'd1230},
{32'd879, 32'd4322, -32'd418, -32'd3480},
{-32'd4833, -32'd7435, 32'd3242, 32'd3734},
{-32'd368, 32'd2173, 32'd8180, -32'd2030},
{32'd1641, -32'd4026, 32'd789, -32'd3016},
{32'd6816, 32'd12978, -32'd5087, -32'd798},
{32'd11053, 32'd2384, 32'd2979, 32'd1187},
{-32'd3664, -32'd281, 32'd726, 32'd5560},
{32'd940, 32'd5032, -32'd10708, -32'd1329},
{32'd584, 32'd5169, -32'd173, 32'd1633},
{-32'd6133, -32'd5692, -32'd10527, -32'd1040},
{32'd1165, -32'd7897, -32'd2431, 32'd6945},
{32'd8417, 32'd8056, -32'd3644, 32'd5664},
{-32'd3838, 32'd9056, -32'd2125, 32'd3988},
{-32'd4980, 32'd3223, 32'd6225, -32'd5828},
{-32'd9505, -32'd5205, -32'd9159, 32'd60},
{32'd6351, 32'd1080, 32'd1870, 32'd1912},
{-32'd3775, 32'd2756, 32'd2724, 32'd5113},
{32'd4860, -32'd6018, 32'd4603, 32'd3864},
{32'd6792, -32'd5400, 32'd2943, 32'd1633},
{-32'd1881, 32'd8080, -32'd16415, -32'd5417}
},
{{32'd8237, -32'd1371, 32'd4995, 32'd214},
{32'd1091, -32'd2281, -32'd3958, -32'd4170},
{-32'd8046, -32'd1558, -32'd1874, 32'd690},
{32'd1, 32'd7142, 32'd7989, 32'd1602},
{-32'd12922, 32'd284, -32'd1572, 32'd584},
{-32'd4241, 32'd2641, 32'd2168, 32'd1514},
{32'd8542, -32'd3050, 32'd1971, 32'd1321},
{32'd1723, -32'd6896, -32'd284, -32'd7319},
{-32'd752, 32'd932, -32'd5040, 32'd5959},
{32'd8608, 32'd6591, 32'd5824, 32'd5592},
{32'd2469, -32'd6187, 32'd591, -32'd1995},
{32'd1741, 32'd8012, 32'd6024, 32'd734},
{32'd794, 32'd4822, 32'd1809, -32'd99},
{-32'd9984, -32'd2736, 32'd993, -32'd3997},
{-32'd6961, -32'd2610, -32'd5014, -32'd1709},
{32'd9301, -32'd7428, -32'd301, -32'd8605},
{32'd7007, -32'd445, 32'd475, 32'd3888},
{32'd13118, 32'd1146, 32'd2655, 32'd3769},
{32'd2600, 32'd3978, -32'd7331, 32'd3102},
{32'd5016, 32'd3647, -32'd3697, 32'd3767},
{-32'd5983, 32'd7219, -32'd717, 32'd3138},
{-32'd1783, -32'd5934, -32'd1335, 32'd4215},
{32'd2125, 32'd891, -32'd12202, -32'd3898},
{32'd2679, -32'd2624, -32'd3578, -32'd714},
{-32'd2178, 32'd3136, 32'd6778, 32'd2011},
{32'd7886, 32'd2454, -32'd1200, -32'd3870},
{32'd3484, -32'd6334, -32'd9370, -32'd219},
{-32'd703, -32'd2715, -32'd5342, -32'd937},
{32'd1916, 32'd4878, 32'd2767, 32'd2459},
{-32'd10955, 32'd5562, 32'd819, 32'd1410},
{32'd7788, 32'd4510, 32'd4467, -32'd6747},
{-32'd6360, -32'd666, -32'd3947, -32'd2354},
{32'd1367, -32'd4040, 32'd7233, 32'd3874},
{-32'd7047, 32'd2011, 32'd3230, -32'd2105},
{32'd6230, 32'd2882, 32'd9863, 32'd6396},
{32'd2318, -32'd3859, -32'd522, 32'd1172},
{-32'd8119, -32'd14004, 32'd1844, -32'd5770},
{-32'd2876, -32'd1146, 32'd9059, 32'd74},
{32'd5039, 32'd5291, 32'd4864, 32'd826},
{32'd3484, 32'd313, -32'd1981, 32'd890},
{-32'd8084, -32'd486, 32'd27, -32'd1366},
{32'd7865, 32'd2249, -32'd1876, 32'd7703},
{32'd9869, 32'd2552, -32'd7683, 32'd6986},
{32'd2116, -32'd2660, -32'd5692, -32'd4310},
{32'd373, -32'd6055, -32'd2793, 32'd311},
{32'd2477, 32'd5697, 32'd998, -32'd139},
{32'd2161, -32'd3205, -32'd9505, -32'd1075},
{32'd2006, 32'd4542, -32'd2396, -32'd577},
{32'd12287, 32'd620, 32'd865, 32'd4600},
{-32'd2804, 32'd39, -32'd3996, 32'd428},
{32'd4209, 32'd1219, -32'd6138, 32'd5239},
{-32'd4935, -32'd2117, 32'd5359, -32'd254},
{32'd4511, -32'd10179, 32'd1124, 32'd3497},
{32'd299, 32'd4348, -32'd2301, 32'd1393},
{-32'd6879, 32'd2955, 32'd4901, 32'd1400},
{-32'd3294, -32'd4249, -32'd4351, -32'd4001},
{32'd887, -32'd3347, 32'd1644, -32'd2421},
{-32'd18642, 32'd1702, -32'd6378, -32'd5364},
{32'd1475, -32'd9991, -32'd5050, -32'd543},
{-32'd3450, 32'd709, -32'd2106, -32'd4046},
{32'd1801, -32'd3028, -32'd4938, 32'd4073},
{-32'd2534, -32'd1848, 32'd2935, 32'd1796},
{-32'd2978, -32'd6401, -32'd11917, -32'd5289},
{-32'd2744, 32'd2642, -32'd5250, 32'd1874},
{32'd8071, 32'd4410, 32'd1994, -32'd3101},
{32'd2028, 32'd9059, 32'd3174, 32'd4176},
{-32'd2946, -32'd628, -32'd1210, -32'd1277},
{32'd2636, -32'd3121, 32'd1404, -32'd1657},
{32'd13397, 32'd415, -32'd1825, -32'd4557},
{-32'd9665, -32'd1267, 32'd3696, 32'd258},
{-32'd17904, -32'd3685, 32'd8737, -32'd2199},
{32'd2499, -32'd3539, 32'd1318, 32'd2773},
{32'd8573, 32'd5863, -32'd298, -32'd3955},
{32'd8095, -32'd1639, -32'd1941, 32'd757},
{-32'd710, -32'd3542, 32'd4133, -32'd1504},
{-32'd2025, -32'd727, -32'd1508, -32'd9352},
{-32'd9654, -32'd8679, -32'd4284, -32'd2308},
{-32'd8545, 32'd2678, -32'd4088, 32'd569},
{-32'd2028, 32'd6450, 32'd9264, -32'd1558},
{32'd1631, -32'd280, 32'd759, 32'd1977},
{32'd3335, 32'd3849, 32'd2338, -32'd1043},
{32'd8669, 32'd11204, -32'd5469, -32'd1758},
{-32'd8130, -32'd240, 32'd1698, -32'd733},
{32'd4019, -32'd2226, 32'd317, 32'd1518},
{-32'd9890, -32'd2068, -32'd845, -32'd199},
{-32'd707, 32'd17646, -32'd2412, 32'd5106},
{32'd3797, 32'd1346, 32'd8840, 32'd7796},
{-32'd7730, -32'd7742, -32'd1633, -32'd4891},
{-32'd102, -32'd281, -32'd1053, -32'd8983},
{32'd7408, 32'd6554, -32'd4456, -32'd1437},
{32'd9073, 32'd2991, 32'd1475, 32'd3858},
{-32'd4135, -32'd1786, -32'd8609, 32'd1198},
{-32'd61, -32'd3286, 32'd3353, 32'd2428},
{-32'd1695, -32'd3189, 32'd4435, 32'd1931},
{32'd13259, -32'd6486, -32'd1912, 32'd2616},
{32'd7447, -32'd2438, -32'd395, -32'd2134},
{32'd7013, 32'd541, 32'd8137, 32'd5223},
{-32'd2935, -32'd8386, 32'd4998, -32'd1534},
{32'd175, 32'd1003, 32'd1348, 32'd3462},
{-32'd2451, 32'd2277, 32'd9048, 32'd3907},
{-32'd1228, -32'd4912, 32'd1707, 32'd1072},
{32'd785, 32'd2264, -32'd6622, 32'd941},
{-32'd7562, 32'd368, -32'd3708, -32'd1632},
{32'd6654, 32'd6530, 32'd5152, 32'd2268},
{32'd3657, 32'd4889, -32'd567, -32'd388},
{-32'd7225, -32'd980, -32'd2838, 32'd6457},
{-32'd3769, -32'd6060, -32'd10165, -32'd2782},
{-32'd9221, 32'd7035, -32'd579, -32'd1156},
{32'd1371, 32'd4319, 32'd5293, 32'd2090},
{-32'd751, -32'd1104, -32'd7149, -32'd1602},
{-32'd9823, -32'd2733, -32'd1390, -32'd4301},
{32'd303, -32'd3382, -32'd1094, 32'd3727},
{32'd2437, 32'd2192, 32'd4274, 32'd2666},
{-32'd5027, -32'd8486, -32'd2138, 32'd2604},
{-32'd7033, -32'd3093, -32'd288, 32'd3103},
{-32'd4821, -32'd2724, -32'd6561, -32'd2815},
{-32'd3307, -32'd3734, 32'd2360, 32'd6585},
{32'd2950, 32'd5331, -32'd2113, 32'd831},
{-32'd16169, -32'd3074, 32'd4110, -32'd864},
{32'd12110, -32'd3336, 32'd5873, 32'd7731},
{32'd10942, 32'd7334, 32'd770, -32'd4961},
{-32'd6900, -32'd3504, 32'd6285, 32'd1713},
{32'd225, -32'd1179, -32'd2038, 32'd2787},
{32'd5572, -32'd3479, -32'd3616, -32'd343},
{-32'd6194, -32'd1436, 32'd2486, 32'd3810},
{32'd5825, -32'd4526, -32'd1378, -32'd2297},
{-32'd1118, 32'd1927, -32'd7173, 32'd2550},
{-32'd5318, 32'd1882, -32'd3832, -32'd6751},
{32'd6369, -32'd1927, -32'd4250, -32'd2719},
{-32'd4094, -32'd2888, 32'd520, -32'd5910},
{32'd1389, -32'd1532, -32'd5589, 32'd2144},
{32'd968, -32'd1177, -32'd253, -32'd7888},
{-32'd5798, -32'd8955, 32'd2253, -32'd5761},
{32'd10708, 32'd10195, 32'd1350, -32'd2624},
{-32'd1656, -32'd497, -32'd536, -32'd4539},
{32'd7024, 32'd1495, -32'd5284, 32'd3631},
{-32'd13560, 32'd386, -32'd6331, 32'd2019},
{-32'd6931, 32'd7871, 32'd438, 32'd7573},
{32'd2020, 32'd7374, -32'd7521, 32'd1721},
{-32'd5814, -32'd997, -32'd7179, -32'd6495},
{32'd12805, -32'd793, 32'd4303, 32'd4341},
{-32'd7860, 32'd1867, 32'd1569, -32'd2550},
{32'd588, 32'd1286, -32'd79, -32'd188},
{-32'd2755, -32'd1411, -32'd6636, -32'd215},
{32'd5936, 32'd9112, 32'd7511, 32'd6300},
{-32'd6402, 32'd3538, -32'd2564, 32'd6547},
{-32'd2326, -32'd3668, -32'd6465, -32'd3553},
{-32'd12607, 32'd5843, -32'd6135, 32'd1204},
{32'd3746, 32'd2105, 32'd5002, 32'd1235},
{32'd7828, -32'd4249, -32'd1636, -32'd5178},
{32'd3077, -32'd5937, -32'd4741, -32'd6797},
{32'd10383, 32'd3322, 32'd901, -32'd1176},
{-32'd4764, -32'd1821, -32'd3233, -32'd1077},
{-32'd4414, -32'd2958, 32'd4955, 32'd1328},
{-32'd5029, -32'd4403, -32'd7089, -32'd4314},
{-32'd5931, -32'd4816, 32'd3049, -32'd4832},
{32'd9323, 32'd5526, -32'd362, 32'd805},
{32'd5941, 32'd1336, 32'd5781, 32'd5242},
{-32'd3966, -32'd1808, -32'd2951, 32'd2310},
{-32'd2483, -32'd3340, -32'd4792, 32'd4716},
{-32'd1514, -32'd11149, -32'd2287, -32'd2112},
{32'd1871, 32'd3934, 32'd6855, -32'd968},
{-32'd17622, 32'd1671, -32'd5189, 32'd4594},
{32'd1614, 32'd7846, 32'd3002, -32'd638},
{32'd2109, 32'd1692, 32'd3678, 32'd1023},
{-32'd4728, 32'd3176, -32'd3758, 32'd423},
{-32'd4182, 32'd1004, 32'd7269, -32'd2276},
{32'd1812, -32'd8707, -32'd4105, -32'd6312},
{-32'd8332, -32'd80, 32'd2512, -32'd2122},
{-32'd4772, -32'd2796, 32'd1184, -32'd2277},
{-32'd6476, -32'd3812, 32'd4025, 32'd3555},
{32'd4172, -32'd7349, 32'd385, -32'd1975},
{32'd16102, 32'd5938, 32'd7320, 32'd2197},
{-32'd1777, 32'd2097, -32'd2145, 32'd1907},
{-32'd1179, 32'd5479, -32'd2920, -32'd1312},
{-32'd694, 32'd5198, 32'd3789, -32'd52},
{32'd4541, 32'd4554, -32'd1708, -32'd912},
{-32'd7764, -32'd10071, -32'd1862, -32'd3411},
{32'd11443, -32'd8105, -32'd752, 32'd176},
{-32'd443, -32'd1017, -32'd2385, -32'd4306},
{32'd114, 32'd3125, -32'd10033, -32'd550},
{32'd1780, 32'd2596, -32'd6669, -32'd4345},
{32'd5507, -32'd2562, 32'd472, -32'd1463},
{-32'd2696, -32'd3517, -32'd130, -32'd2842},
{32'd2437, -32'd5510, 32'd1661, -32'd2894},
{-32'd10542, 32'd6051, 32'd4517, 32'd600},
{32'd239, 32'd1176, 32'd1816, 32'd423},
{-32'd9493, -32'd3045, -32'd178, -32'd890},
{32'd942, 32'd4338, -32'd1809, -32'd3032},
{-32'd8063, -32'd4738, -32'd7793, -32'd7505},
{-32'd3946, 32'd1984, -32'd5181, 32'd1464},
{-32'd7617, 32'd3871, -32'd978, -32'd649},
{-32'd9027, 32'd1267, -32'd4980, 32'd1531},
{32'd2170, 32'd5502, 32'd1311, 32'd2827},
{32'd6896, 32'd1651, 32'd651, -32'd2584},
{-32'd6676, 32'd626, 32'd5096, 32'd2534},
{32'd3319, 32'd2118, 32'd2070, -32'd4142},
{32'd10583, 32'd6824, 32'd3615, -32'd140},
{-32'd2126, 32'd137, 32'd7135, -32'd52},
{-32'd1242, -32'd6282, -32'd1739, 32'd2362},
{-32'd8141, -32'd11828, -32'd6301, -32'd6499},
{-32'd1093, -32'd5485, -32'd492, 32'd4866},
{-32'd285, 32'd926, 32'd2883, -32'd2255},
{32'd869, -32'd3447, 32'd8760, 32'd1336},
{32'd10838, 32'd2073, -32'd10823, -32'd144},
{32'd505, 32'd2827, 32'd6594, -32'd3636},
{-32'd9200, -32'd5198, 32'd5303, 32'd2022},
{32'd4089, -32'd3750, 32'd22, -32'd2518},
{-32'd1350, -32'd6106, 32'd1689, -32'd1773},
{32'd5596, -32'd1610, 32'd3551, 32'd709},
{-32'd711, -32'd40, 32'd3741, -32'd2442},
{32'd991, -32'd3161, 32'd210, 32'd1358},
{-32'd14462, 32'd5083, -32'd4148, -32'd3631},
{-32'd8925, -32'd1107, 32'd13940, -32'd705},
{-32'd1515, -32'd2325, -32'd6576, -32'd1648},
{-32'd9112, 32'd3986, -32'd2363, 32'd5187},
{-32'd11987, 32'd306, 32'd2599, -32'd2813},
{32'd33, 32'd7314, -32'd706, -32'd3500},
{32'd7137, 32'd495, 32'd8722, 32'd4273},
{32'd5286, 32'd3965, -32'd3238, 32'd5532},
{-32'd4834, -32'd1833, -32'd1734, -32'd4806},
{-32'd994, -32'd179, -32'd5378, -32'd463},
{32'd5726, -32'd2925, 32'd548, 32'd811},
{-32'd6263, 32'd2961, -32'd6623, -32'd3683},
{32'd12006, -32'd968, -32'd4660, -32'd391},
{32'd7911, 32'd1438, 32'd2380, 32'd1286},
{-32'd2291, 32'd8863, -32'd8507, 32'd728},
{32'd2834, 32'd5013, -32'd4487, -32'd1990},
{32'd796, 32'd5402, 32'd2132, 32'd3168},
{32'd16970, -32'd4797, -32'd1668, 32'd6518},
{-32'd8219, -32'd12339, 32'd703, 32'd1817},
{-32'd11902, 32'd4622, -32'd4267, 32'd713},
{32'd3518, 32'd4733, 32'd1610, -32'd1498},
{-32'd1173, -32'd9586, -32'd6954, 32'd2074},
{32'd4617, -32'd5010, -32'd8635, -32'd7806},
{-32'd7950, -32'd6091, -32'd1316, -32'd4060},
{32'd1365, -32'd1262, 32'd353, -32'd364},
{32'd5367, 32'd2009, 32'd608, 32'd1535},
{32'd5068, 32'd5076, 32'd5863, -32'd226},
{-32'd6415, -32'd899, -32'd12323, 32'd2467},
{-32'd5221, -32'd8107, -32'd789, -32'd679},
{-32'd1917, -32'd8148, -32'd1848, 32'd3296},
{-32'd1457, -32'd4241, -32'd4559, -32'd6089},
{32'd7201, -32'd6569, 32'd3749, -32'd1628},
{32'd4821, 32'd2564, 32'd5284, 32'd2318},
{-32'd4408, -32'd4902, 32'd7068, -32'd6741},
{-32'd9673, -32'd9802, -32'd3281, 32'd114},
{-32'd2260, 32'd10155, -32'd4024, 32'd2667},
{-32'd814, 32'd2424, 32'd7697, 32'd5133},
{32'd11527, 32'd8856, 32'd4839, -32'd372},
{-32'd7725, -32'd776, -32'd9204, 32'd1202},
{32'd1148, 32'd879, -32'd4633, 32'd1796},
{-32'd1558, -32'd747, -32'd1154, -32'd2460},
{-32'd3228, -32'd3425, 32'd1352, 32'd4096},
{-32'd5499, 32'd1380, -32'd6113, -32'd1069},
{-32'd14462, 32'd4227, 32'd381, 32'd1937},
{32'd1588, 32'd5224, -32'd1009, 32'd242},
{32'd4927, 32'd4966, 32'd214, -32'd601},
{-32'd5762, -32'd10192, -32'd4900, -32'd4317},
{32'd3593, -32'd10109, 32'd7673, 32'd1345},
{-32'd714, 32'd2242, 32'd7260, -32'd2149},
{-32'd6218, 32'd3560, -32'd571, 32'd2505},
{32'd214, 32'd1250, -32'd2520, 32'd272},
{32'd720, -32'd2261, 32'd2438, -32'd2271},
{-32'd1360, 32'd3701, -32'd472, -32'd3254},
{32'd5413, 32'd7819, -32'd1788, 32'd9809},
{32'd4596, 32'd2054, 32'd2046, -32'd333},
{-32'd7890, -32'd4388, -32'd678, -32'd117},
{-32'd816, 32'd1883, -32'd78, -32'd5421},
{-32'd3181, -32'd7517, -32'd7206, 32'd6906},
{32'd5462, 32'd9931, -32'd1451, -32'd1975},
{32'd6215, 32'd10129, 32'd1636, -32'd1084},
{32'd4733, 32'd4638, -32'd1281, 32'd1352},
{-32'd10322, -32'd3511, 32'd954, -32'd964},
{32'd3513, 32'd302, -32'd5363, 32'd1173},
{-32'd4068, 32'd3612, -32'd6598, 32'd1798},
{32'd10886, 32'd7933, 32'd8382, 32'd7674},
{32'd5831, -32'd5468, 32'd1797, 32'd3555},
{-32'd280, -32'd1449, -32'd2650, -32'd5074},
{32'd8796, -32'd962, -32'd637, -32'd795},
{32'd4534, 32'd6966, -32'd1130, 32'd6882},
{32'd1814, -32'd2968, -32'd6866, -32'd5760},
{32'd3677, 32'd1136, 32'd473, -32'd2621},
{32'd11072, 32'd8325, -32'd459, 32'd6877},
{32'd4404, 32'd4853, 32'd1738, 32'd2565},
{32'd6165, -32'd4666, -32'd1747, -32'd2732},
{32'd4707, -32'd4238, 32'd2346, -32'd66},
{-32'd5374, -32'd4135, -32'd3401, 32'd4875},
{32'd3669, -32'd1102, -32'd1931, 32'd3749},
{-32'd4020, -32'd1505, 32'd2381, -32'd864},
{-32'd5238, -32'd8698, -32'd2774, -32'd1734},
{32'd5288, 32'd4029, 32'd3420, 32'd3376},
{32'd8514, 32'd11007, -32'd4728, 32'd118},
{-32'd5716, -32'd2396, -32'd2232, -32'd164},
{-32'd518, 32'd4439, -32'd1309, 32'd3261},
{-32'd3372, -32'd6467, 32'd4050, -32'd1517},
{-32'd4867, -32'd5173, 32'd1485, -32'd2486},
{-32'd1492, -32'd1298, 32'd11525, 32'd6385},
{32'd5427, 32'd3173, 32'd10895, 32'd5642},
{-32'd967, -32'd3205, -32'd3630, 32'd50}
},
{{32'd6498, 32'd6622, -32'd4281, 32'd7305},
{-32'd4268, 32'd1137, -32'd6473, 32'd915},
{32'd4004, -32'd5565, -32'd267, -32'd2112},
{32'd11429, 32'd6151, -32'd1670, 32'd6686},
{-32'd934, -32'd1364, 32'd885, 32'd2436},
{-32'd3452, -32'd1303, -32'd2127, 32'd6493},
{-32'd1079, -32'd181, 32'd8593, 32'd1345},
{-32'd10625, -32'd9851, 32'd11147, 32'd4720},
{32'd6427, -32'd2239, -32'd5714, -32'd7280},
{32'd6507, 32'd11912, 32'd3454, 32'd10612},
{-32'd19978, 32'd1193, 32'd6691, -32'd539},
{-32'd3295, -32'd9085, 32'd4585, -32'd6260},
{32'd2636, 32'd3617, -32'd7370, -32'd2988},
{-32'd4069, -32'd4424, -32'd8760, -32'd2380},
{-32'd6934, 32'd375, -32'd9033, -32'd1368},
{32'd6394, 32'd3923, -32'd882, -32'd16202},
{32'd6854, -32'd429, -32'd4331, -32'd3865},
{32'd3814, -32'd3867, 32'd773, 32'd1752},
{32'd2435, 32'd3309, 32'd4212, 32'd7205},
{-32'd24003, -32'd4533, 32'd437, 32'd6511},
{32'd72, -32'd1876, 32'd1468, 32'd13514},
{-32'd13374, -32'd7547, -32'd6651, -32'd3825},
{32'd1415, -32'd6415, -32'd7586, -32'd2196},
{32'd4291, 32'd7070, 32'd4482, 32'd3697},
{32'd2716, 32'd4317, 32'd7728, 32'd2273},
{-32'd3700, 32'd8692, -32'd3565, 32'd123},
{-32'd2751, -32'd4356, 32'd6737, 32'd3731},
{32'd11594, -32'd2074, 32'd11783, 32'd5687},
{-32'd3610, -32'd2598, 32'd4801, 32'd4539},
{-32'd651, 32'd449, 32'd945, -32'd1005},
{32'd1656, -32'd12781, -32'd14387, -32'd2332},
{-32'd12676, -32'd9697, -32'd2907, -32'd5169},
{32'd4982, 32'd14417, 32'd14586, 32'd788},
{-32'd949, -32'd4801, -32'd1701, -32'd9185},
{-32'd2493, 32'd6611, 32'd5899, 32'd688},
{-32'd15723, -32'd15258, 32'd1042, 32'd5929},
{32'd3963, -32'd1335, 32'd9772, 32'd2695},
{-32'd2534, -32'd749, -32'd3671, -32'd4451},
{-32'd1603, 32'd11824, 32'd7522, 32'd1609},
{32'd5142, 32'd11021, 32'd3004, -32'd1427},
{-32'd3696, 32'd1501, -32'd281, 32'd5372},
{-32'd13090, 32'd7127, 32'd4135, -32'd817},
{-32'd3419, 32'd6961, 32'd5349, -32'd2263},
{32'd7340, -32'd4774, -32'd3336, -32'd1816},
{32'd2492, -32'd4196, -32'd8392, -32'd5114},
{-32'd7692, 32'd1345, -32'd9390, -32'd3746},
{-32'd11685, -32'd5044, 32'd1357, 32'd10631},
{-32'd4359, 32'd3048, -32'd4582, -32'd6812},
{-32'd10423, 32'd11328, 32'd3262, 32'd4308},
{-32'd12119, -32'd9212, -32'd5444, 32'd1759},
{-32'd5221, -32'd6510, -32'd11099, -32'd3376},
{32'd3543, -32'd465, 32'd6103, -32'd1506},
{32'd3907, -32'd3612, -32'd4466, -32'd9888},
{32'd8521, 32'd11641, 32'd5073, 32'd4670},
{32'd4937, -32'd9190, 32'd243, 32'd12726},
{-32'd8114, 32'd7373, -32'd7337, -32'd3884},
{-32'd8, 32'd2069, -32'd367, 32'd3422},
{-32'd1126, 32'd1126, -32'd935, -32'd6899},
{32'd2853, 32'd8007, -32'd9783, -32'd2766},
{-32'd3528, 32'd1735, -32'd4475, -32'd3690},
{-32'd1972, -32'd10775, 32'd4172, 32'd5961},
{32'd10949, -32'd353, 32'd635, -32'd2150},
{-32'd16999, -32'd7023, -32'd1215, -32'd7455},
{-32'd4389, -32'd1892, -32'd12521, 32'd7975},
{-32'd1656, 32'd7442, -32'd10789, 32'd1630},
{-32'd1934, 32'd9942, 32'd8674, 32'd1711},
{-32'd6266, -32'd9105, -32'd5022, 32'd12172},
{-32'd900, -32'd5767, 32'd940, -32'd1699},
{-32'd3004, -32'd4607, 32'd1678, 32'd1286},
{32'd10, -32'd4607, 32'd9896, 32'd3764},
{-32'd1572, 32'd7215, 32'd8505, 32'd242},
{-32'd5000, 32'd1506, 32'd14, 32'd345},
{32'd1161, -32'd6470, -32'd1131, -32'd6312},
{-32'd1766, -32'd100, 32'd2338, 32'd434},
{-32'd1837, -32'd1115, -32'd2568, -32'd1706},
{32'd3765, 32'd12256, -32'd15825, -32'd11101},
{32'd2631, -32'd9275, 32'd8317, 32'd1692},
{-32'd2750, -32'd861, -32'd2893, -32'd10333},
{32'd17042, 32'd6425, 32'd11229, 32'd8527},
{-32'd9929, -32'd2975, -32'd4925, -32'd1425},
{32'd12013, 32'd3541, 32'd8422, 32'd8514},
{32'd10503, 32'd15081, 32'd5451, -32'd5169},
{-32'd7456, 32'd154, 32'd3831, 32'd10110},
{32'd3167, -32'd376, 32'd1902, -32'd9756},
{32'd5258, -32'd4557, -32'd2681, -32'd7168},
{-32'd18747, -32'd4360, -32'd10360, 32'd498},
{-32'd16929, 32'd5832, -32'd5605, 32'd6742},
{32'd2207, 32'd3313, 32'd2615, 32'd4461},
{32'd1429, -32'd3511, -32'd3404, 32'd4569},
{32'd11918, -32'd11508, 32'd6050, -32'd5991},
{32'd9908, 32'd5086, -32'd5555, -32'd297},
{-32'd1937, -32'd2253, 32'd2603, -32'd2470},
{-32'd2138, -32'd7020, -32'd7801, -32'd13312},
{-32'd2577, 32'd4861, 32'd6250, -32'd4685},
{32'd6578, -32'd3429, 32'd856, 32'd1794},
{-32'd668, -32'd2334, 32'd7796, -32'd4298},
{32'd8176, 32'd2829, -32'd2953, -32'd1583},
{32'd10271, -32'd387, -32'd1976, 32'd639},
{-32'd3210, 32'd606, 32'd10626, -32'd9283},
{32'd7665, 32'd2481, -32'd4000, -32'd6065},
{-32'd2813, 32'd5891, -32'd8999, 32'd6510},
{-32'd6665, -32'd3764, -32'd5553, -32'd4210},
{32'd17829, 32'd13838, 32'd2851, 32'd19378},
{-32'd449, 32'd2108, -32'd385, 32'd8795},
{-32'd3640, 32'd5287, 32'd8464, 32'd3662},
{-32'd4125, 32'd627, -32'd714, 32'd1733},
{-32'd12504, -32'd10728, -32'd766, 32'd6209},
{-32'd12908, -32'd13575, 32'd5019, -32'd4526},
{-32'd1510, 32'd11161, 32'd4090, 32'd3494},
{-32'd7115, -32'd7307, -32'd8932, -32'd4038},
{32'd4276, 32'd4219, 32'd13183, -32'd8650},
{32'd1268, 32'd11539, 32'd8898, 32'd5091},
{32'd7193, 32'd12443, -32'd3863, 32'd15477},
{32'd1559, 32'd6194, 32'd2128, 32'd4489},
{-32'd4352, 32'd2830, -32'd152, 32'd5249},
{32'd3118, -32'd1058, -32'd2774, -32'd7885},
{-32'd607, -32'd4130, -32'd9304, -32'd4407},
{-32'd5847, -32'd12960, -32'd1132, -32'd5803},
{32'd3657, 32'd3509, 32'd946, -32'd875},
{32'd3842, 32'd3583, -32'd2988, -32'd4291},
{-32'd5698, -32'd899, 32'd547, -32'd2189},
{32'd13256, 32'd1195, -32'd509, -32'd7105},
{-32'd1556, -32'd13333, 32'd3509, -32'd1507},
{-32'd781, -32'd4251, -32'd6479, 32'd1481},
{-32'd11878, 32'd1188, 32'd8028, 32'd5170},
{32'd16657, 32'd618, -32'd9418, 32'd9511},
{-32'd818, 32'd10897, -32'd5602, -32'd6039},
{-32'd7944, -32'd3780, -32'd2941, -32'd7477},
{32'd5968, -32'd8497, 32'd288, -32'd2960},
{32'd4036, 32'd4516, -32'd3128, -32'd2145},
{-32'd12524, -32'd16671, -32'd1213, -32'd7967},
{-32'd9166, 32'd1334, 32'd7414, 32'd1373},
{32'd435, -32'd3797, -32'd3259, 32'd319},
{32'd1010, 32'd1977, 32'd14683, 32'd4850},
{32'd4530, 32'd976, -32'd5168, 32'd1089},
{-32'd577, 32'd9716, 32'd5078, -32'd2330},
{-32'd8888, -32'd7990, 32'd1951, 32'd5793},
{32'd10342, -32'd3077, -32'd7947, 32'd665},
{-32'd3902, -32'd14797, 32'd4387, -32'd9376},
{-32'd20988, -32'd3619, 32'd5361, 32'd2471},
{-32'd6984, 32'd10113, 32'd13737, -32'd12886},
{32'd4336, 32'd4155, 32'd12793, 32'd3917},
{-32'd5757, 32'd186, -32'd3238, -32'd4878},
{-32'd13441, -32'd5243, 32'd5390, -32'd4786},
{32'd14268, 32'd10553, 32'd1769, 32'd7525},
{32'd9477, 32'd329, -32'd481, -32'd11319},
{-32'd6244, -32'd715, -32'd8479, -32'd5666},
{-32'd2322, -32'd9308, -32'd8227, -32'd4581},
{32'd13643, -32'd2126, 32'd9610, 32'd7624},
{-32'd365, -32'd15792, -32'd2712, 32'd410},
{32'd3274, -32'd4561, 32'd1472, -32'd5803},
{32'd8753, -32'd2734, 32'd9469, 32'd735},
{32'd3406, 32'd3555, 32'd5575, -32'd11859},
{-32'd11244, -32'd1674, -32'd12292, -32'd1010},
{-32'd13872, -32'd3191, -32'd7459, -32'd8314},
{32'd4888, 32'd1078, -32'd848, 32'd5536},
{-32'd6990, 32'd399, 32'd11058, 32'd2693},
{-32'd4, -32'd3134, 32'd9593, 32'd9093},
{32'd7098, -32'd5435, -32'd8507, -32'd5952},
{-32'd6202, 32'd5117, -32'd8005, -32'd8303},
{-32'd19245, -32'd5741, 32'd4472, 32'd1884},
{32'd21056, -32'd1274, -32'd2060, -32'd5915},
{-32'd14934, 32'd1308, -32'd2190, 32'd4176},
{32'd15567, 32'd3473, 32'd6987, 32'd15950},
{-32'd10129, -32'd8514, 32'd6509, 32'd1936},
{-32'd7099, -32'd8118, 32'd8805, 32'd1636},
{-32'd1737, -32'd6616, 32'd6181, 32'd292},
{-32'd7233, 32'd127, -32'd225, -32'd5821},
{32'd13334, 32'd15474, -32'd16597, -32'd3671},
{-32'd7890, -32'd16255, -32'd6274, -32'd337},
{-32'd2526, -32'd14444, 32'd1490, -32'd10596},
{-32'd7859, -32'd2850, 32'd20397, 32'd7083},
{32'd6738, 32'd7094, 32'd2054, 32'd6630},
{32'd10735, -32'd1841, 32'd201, 32'd6043},
{32'd3994, 32'd3683, 32'd2764, 32'd13151},
{-32'd746, 32'd2384, -32'd11817, -32'd3397},
{32'd10928, 32'd7489, 32'd6809, 32'd7429},
{32'd2466, -32'd11886, 32'd2593, -32'd2865},
{32'd180, 32'd736, -32'd9068, 32'd2886},
{-32'd428, -32'd5239, 32'd1844, -32'd4945},
{32'd15209, 32'd13679, 32'd8527, -32'd3198},
{-32'd3430, -32'd3597, -32'd6012, -32'd7271},
{-32'd1210, 32'd4449, -32'd1772, 32'd9707},
{-32'd2012, 32'd15326, -32'd12442, -32'd2679},
{32'd7100, -32'd4323, 32'd4318, -32'd1111},
{32'd9409, -32'd9945, 32'd608, -32'd1656},
{-32'd5507, -32'd4002, -32'd7271, 32'd3351},
{32'd1369, -32'd7466, -32'd6010, -32'd435},
{32'd11079, 32'd4491, 32'd3193, 32'd1312},
{-32'd4365, 32'd3052, -32'd7533, 32'd14096},
{32'd8870, -32'd6689, 32'd6123, -32'd745},
{32'd4074, -32'd630, 32'd5799, -32'd1631},
{32'd4135, -32'd1437, -32'd7948, -32'd2697},
{-32'd507, -32'd4665, -32'd5722, 32'd4645},
{32'd5208, -32'd4393, -32'd1773, -32'd2595},
{-32'd5160, -32'd1847, 32'd6447, 32'd1043},
{-32'd1814, 32'd1851, -32'd4508, -32'd1413},
{-32'd602, -32'd3727, 32'd5303, 32'd1571},
{-32'd5325, 32'd1618, 32'd1673, 32'd1296},
{-32'd283, -32'd497, 32'd1997, -32'd3343},
{-32'd10554, -32'd1725, -32'd6881, -32'd3389},
{32'd5249, 32'd1179, -32'd3061, -32'd6993},
{32'd3699, 32'd1437, 32'd7129, -32'd10886},
{-32'd13688, 32'd2912, 32'd6495, 32'd15035},
{32'd5065, -32'd283, 32'd7216, -32'd1906},
{-32'd25597, 32'd8463, 32'd1501, 32'd5352},
{-32'd635, -32'd3552, -32'd4339, -32'd5893},
{32'd3632, -32'd3758, -32'd5604, 32'd2220},
{32'd6521, -32'd1586, 32'd7215, 32'd2202},
{32'd1170, 32'd2951, -32'd907, -32'd3168},
{-32'd4864, 32'd2032, -32'd1767, -32'd10836},
{-32'd8848, 32'd2084, -32'd3937, 32'd263},
{-32'd15457, 32'd694, 32'd9729, 32'd2690},
{-32'd2255, -32'd6045, 32'd3462, -32'd913},
{32'd587, 32'd4785, -32'd313, -32'd5649},
{-32'd4027, -32'd11445, -32'd5635, 32'd9579},
{32'd3726, 32'd7059, 32'd1001, 32'd14603},
{-32'd3485, -32'd9805, 32'd12481, -32'd9474},
{-32'd817, -32'd1342, -32'd8868, 32'd9724},
{32'd2295, -32'd12521, 32'd116, -32'd5270},
{-32'd6387, -32'd4694, -32'd13884, 32'd3351},
{-32'd8312, 32'd5725, 32'd4180, 32'd6491},
{32'd10561, 32'd2341, 32'd9495, 32'd4647},
{32'd2602, -32'd18274, 32'd5144, -32'd3227},
{-32'd970, -32'd14237, -32'd8074, 32'd8683},
{32'd2351, 32'd4456, 32'd7930, 32'd9115},
{-32'd9618, 32'd201, -32'd6800, -32'd4779},
{-32'd605, 32'd4012, -32'd3356, -32'd5402},
{-32'd5068, 32'd3345, 32'd16462, 32'd3211},
{-32'd5202, 32'd1697, -32'd9830, -32'd5052},
{-32'd20543, -32'd14953, 32'd4941, 32'd756},
{-32'd3163, 32'd2463, 32'd9613, -32'd11163},
{32'd2349, 32'd7400, -32'd760, -32'd1549},
{-32'd971, -32'd505, 32'd3132, -32'd5565},
{32'd6961, -32'd6266, 32'd7250, -32'd4000},
{-32'd10124, -32'd5535, -32'd18110, -32'd470},
{-32'd87, -32'd9261, 32'd2829, 32'd7363},
{-32'd1707, 32'd4668, 32'd12130, 32'd12399},
{32'd12728, 32'd956, -32'd1554, 32'd2046},
{32'd22262, 32'd10008, -32'd8582, -32'd12564},
{-32'd8989, 32'd5566, 32'd13057, 32'd2592},
{-32'd7041, 32'd1938, -32'd13753, 32'd1999},
{32'd6270, -32'd4056, -32'd6014, -32'd1033},
{32'd10441, 32'd4305, -32'd9321, -32'd7682},
{32'd2315, 32'd14924, 32'd6969, 32'd9545},
{32'd9665, 32'd7039, 32'd4946, 32'd7710},
{-32'd3000, -32'd6807, 32'd3117, 32'd2276},
{-32'd7193, -32'd6328, -32'd3642, 32'd1},
{-32'd6831, 32'd2560, 32'd3967, 32'd14621},
{32'd737, 32'd4952, -32'd9408, 32'd7220},
{32'd1182, 32'd2063, -32'd6084, -32'd5339},
{-32'd2686, -32'd2691, 32'd2022, 32'd3733},
{32'd11457, -32'd5828, -32'd582, -32'd2942},
{-32'd2440, 32'd9578, 32'd11678, 32'd15780},
{-32'd13102, 32'd2152, 32'd2436, -32'd12343},
{-32'd9867, -32'd1128, -32'd2148, 32'd17634},
{32'd6341, 32'd163, 32'd6241, 32'd1558},
{32'd8935, 32'd1668, -32'd201, -32'd2746},
{-32'd7909, 32'd818, 32'd11460, -32'd2586},
{32'd5076, -32'd250, -32'd11330, -32'd1711},
{-32'd10029, -32'd11428, -32'd4293, -32'd513},
{32'd11720, 32'd5929, -32'd4058, 32'd3406},
{-32'd3635, -32'd3823, 32'd1077, -32'd8682},
{-32'd642, 32'd3329, 32'd10298, -32'd4956},
{32'd18911, -32'd5955, 32'd8916, -32'd10809},
{32'd7660, -32'd1425, -32'd4617, -32'd3144},
{32'd8293, 32'd6794, 32'd9964, 32'd824},
{-32'd575, 32'd7709, 32'd2520, -32'd13042},
{-32'd15456, -32'd6067, -32'd2650, -32'd8900},
{-32'd1149, 32'd3602, -32'd7269, 32'd1837},
{32'd6288, -32'd6283, 32'd11094, 32'd3343},
{32'd3033, -32'd4084, 32'd6666, -32'd3843},
{-32'd6950, -32'd9324, -32'd2880, 32'd5407},
{32'd8678, -32'd255, -32'd4842, -32'd14804},
{32'd12597, 32'd1858, 32'd3370, 32'd121},
{-32'd5881, -32'd269, 32'd9631, 32'd2927},
{32'd6600, 32'd13716, 32'd5156, 32'd4433},
{-32'd2234, -32'd16043, 32'd1364, -32'd781},
{32'd5463, -32'd7523, 32'd455, -32'd7825},
{32'd1242, -32'd5034, -32'd3512, -32'd8236},
{-32'd68, -32'd2322, 32'd3353, 32'd4400},
{-32'd13289, -32'd1635, 32'd8243, 32'd1581},
{-32'd1578, 32'd1429, 32'd6158, -32'd10282},
{32'd6213, 32'd308, -32'd4465, 32'd5503},
{-32'd707, 32'd3952, 32'd7405, -32'd6321},
{32'd8565, 32'd3799, -32'd2965, -32'd9149},
{32'd11025, -32'd3400, 32'd6972, -32'd9112},
{-32'd5277, 32'd867, 32'd4171, -32'd4966},
{32'd8335, 32'd11302, -32'd385, 32'd3475},
{-32'd4407, -32'd459, -32'd1399, 32'd5188},
{32'd7209, 32'd1413, -32'd4262, 32'd2691},
{32'd10325, 32'd16947, 32'd7959, 32'd10460},
{-32'd873, -32'd1914, -32'd1100, -32'd2818},
{-32'd2915, -32'd1367, -32'd3903, 32'd6100},
{32'd6015, -32'd476, -32'd1653, -32'd5882},
{-32'd762, 32'd4270, 32'd2717, -32'd5137},
{-32'd55, -32'd9480, 32'd134, -32'd9797},
{-32'd9801, 32'd7714, 32'd3246, 32'd3504},
{32'd3103, -32'd8136, 32'd1204, 32'd3985},
{32'd5870, 32'd9298, 32'd5332, 32'd77}
},
{{32'd9485, 32'd12332, 32'd5113, 32'd4015},
{32'd3720, -32'd5305, -32'd7796, -32'd10142},
{32'd1917, -32'd58, -32'd4630, -32'd5437},
{32'd3627, 32'd178, 32'd14214, 32'd286},
{32'd5133, -32'd15574, -32'd10201, -32'd4828},
{32'd549, 32'd5484, -32'd14946, -32'd6811},
{32'd303, 32'd9787, 32'd322, 32'd10199},
{-32'd6462, 32'd14921, 32'd8182, 32'd6881},
{-32'd5792, -32'd3186, -32'd972, 32'd3756},
{32'd7593, -32'd1788, 32'd108, 32'd5403},
{-32'd4397, 32'd2798, -32'd13616, 32'd8491},
{-32'd10212, 32'd7478, 32'd202, 32'd2024},
{-32'd12681, -32'd2995, 32'd8566, -32'd11331},
{-32'd3137, -32'd15104, 32'd4033, 32'd1972},
{-32'd14413, -32'd5692, 32'd4827, -32'd3738},
{32'd4554, 32'd2470, 32'd4888, 32'd402},
{32'd2578, 32'd4960, 32'd4123, -32'd7866},
{-32'd12993, -32'd4087, 32'd20506, -32'd8851},
{32'd1789, -32'd19490, 32'd12341, 32'd6318},
{-32'd4629, -32'd2443, -32'd6409, 32'd753},
{-32'd4873, -32'd6844, 32'd146, 32'd1164},
{-32'd1581, 32'd8419, 32'd907, -32'd9699},
{32'd8553, 32'd4065, 32'd103, -32'd277},
{-32'd2182, 32'd5127, -32'd963, -32'd2655},
{32'd1150, 32'd7725, 32'd5869, 32'd3073},
{32'd820, 32'd7941, 32'd6614, 32'd5409},
{-32'd12317, -32'd9780, -32'd3757, 32'd9667},
{-32'd806, 32'd9539, 32'd5771, 32'd711},
{-32'd178, -32'd1765, 32'd1358, -32'd7705},
{-32'd411, -32'd499, 32'd6745, -32'd310},
{-32'd3080, -32'd4136, 32'd8598, 32'd468},
{-32'd8916, -32'd2864, 32'd9030, -32'd8484},
{32'd10302, 32'd8742, 32'd645, 32'd15742},
{-32'd5437, 32'd9156, -32'd7415, -32'd214},
{-32'd8380, 32'd5164, 32'd7093, -32'd2008},
{32'd9407, 32'd1121, 32'd11505, -32'd14723},
{-32'd4508, 32'd2738, -32'd4156, 32'd12677},
{32'd10780, -32'd8042, -32'd5114, -32'd4555},
{-32'd2694, -32'd3882, -32'd6724, -32'd4880},
{32'd3148, 32'd4817, -32'd8121, 32'd4625},
{32'd7492, -32'd10147, -32'd3460, -32'd9},
{32'd3657, -32'd3507, 32'd11497, 32'd3876},
{-32'd306, -32'd5350, -32'd5069, -32'd5078},
{-32'd3653, 32'd4175, -32'd2573, 32'd2355},
{-32'd14503, -32'd10267, -32'd10596, -32'd790},
{32'd2272, -32'd16345, -32'd11553, 32'd3426},
{-32'd14919, -32'd343, -32'd7047, -32'd5323},
{-32'd6390, -32'd11931, 32'd8402, -32'd1276},
{-32'd12284, -32'd2415, -32'd5903, -32'd8423},
{-32'd87, -32'd2334, 32'd8929, 32'd2379},
{-32'd16419, -32'd1349, 32'd8749, -32'd1301},
{-32'd19, 32'd2807, 32'd6082, -32'd3042},
{-32'd8835, 32'd4431, 32'd2954, -32'd409},
{-32'd251, 32'd1825, 32'd8209, -32'd8456},
{32'd1248, 32'd1621, 32'd9705, -32'd214},
{32'd15651, -32'd7254, 32'd1193, 32'd5704},
{32'd488, 32'd4774, -32'd190, -32'd1309},
{-32'd5327, -32'd7744, 32'd15497, -32'd848},
{32'd1793, -32'd8374, 32'd2152, 32'd8800},
{32'd2446, -32'd7807, -32'd11860, -32'd5543},
{32'd5379, -32'd2566, 32'd14218, 32'd1043},
{-32'd640, 32'd6555, 32'd6579, -32'd3814},
{-32'd12187, -32'd12046, 32'd98, -32'd12755},
{-32'd438, -32'd7147, -32'd2881, -32'd7434},
{-32'd10549, 32'd15853, -32'd303, -32'd2480},
{-32'd7428, 32'd20724, 32'd10320, -32'd5046},
{32'd2441, -32'd7743, -32'd16690, 32'd11144},
{-32'd10321, 32'd13373, -32'd10566, -32'd6912},
{-32'd1010, 32'd11130, 32'd2169, -32'd1931},
{-32'd11139, 32'd16695, 32'd9107, 32'd11361},
{32'd15579, 32'd1172, -32'd926, 32'd5457},
{32'd4343, 32'd4319, 32'd3678, 32'd4110},
{-32'd5716, -32'd1760, 32'd2671, -32'd3445},
{32'd8228, 32'd1849, -32'd35, 32'd4385},
{32'd679, 32'd7022, -32'd701, 32'd5279},
{32'd5280, -32'd3791, 32'd5398, -32'd7481},
{-32'd9342, -32'd4707, -32'd1293, -32'd6499},
{32'd2424, -32'd9557, -32'd7036, -32'd6145},
{-32'd3038, 32'd4998, 32'd6083, 32'd4140},
{-32'd6943, 32'd773, 32'd1268, 32'd4874},
{32'd3606, -32'd6875, -32'd2622, 32'd2562},
{32'd10598, -32'd15165, 32'd4391, -32'd2899},
{-32'd4129, -32'd7125, -32'd6683, 32'd6562},
{-32'd1006, 32'd4559, 32'd5734, -32'd3752},
{-32'd3602, -32'd3699, 32'd2970, -32'd5511},
{32'd1825, -32'd15121, 32'd17271, 32'd488},
{-32'd3564, 32'd3657, 32'd14265, -32'd900},
{-32'd12535, -32'd10395, 32'd6583, -32'd12386},
{-32'd17901, -32'd9464, -32'd2229, -32'd5323},
{32'd13, -32'd6335, 32'd6020, -32'd459},
{32'd3431, 32'd1673, -32'd8811, 32'd2225},
{32'd14374, -32'd605, -32'd4450, -32'd19916},
{-32'd5224, -32'd3254, -32'd2706, -32'd4135},
{32'd3286, 32'd15847, 32'd467, -32'd6097},
{-32'd6946, -32'd3597, 32'd2970, -32'd10790},
{32'd1373, 32'd3372, -32'd7989, 32'd794},
{32'd5950, -32'd2723, -32'd7079, -32'd2536},
{-32'd3291, 32'd10585, 32'd197, 32'd2796},
{-32'd7507, 32'd4723, 32'd4022, -32'd13372},
{32'd319, -32'd3757, -32'd7262, 32'd3904},
{-32'd3735, 32'd159, -32'd2840, -32'd566},
{-32'd1440, 32'd7026, 32'd5389, -32'd3728},
{32'd1597, 32'd5094, -32'd11337, 32'd10401},
{-32'd5008, -32'd420, 32'd3834, -32'd3062},
{32'd839, 32'd2551, 32'd2017, 32'd16838},
{32'd11586, -32'd2832, -32'd5700, 32'd3211},
{32'd1687, -32'd19691, 32'd1744, 32'd3516},
{32'd11655, -32'd3014, -32'd5303, 32'd4226},
{-32'd3809, -32'd6478, -32'd12951, 32'd9260},
{32'd2773, 32'd8706, -32'd1316, -32'd5503},
{-32'd3321, -32'd10879, 32'd1769, 32'd5565},
{-32'd5836, -32'd7399, -32'd2905, 32'd2869},
{32'd11643, 32'd10676, -32'd2665, 32'd6229},
{32'd4735, -32'd1785, -32'd6458, -32'd9428},
{-32'd2126, -32'd18424, 32'd5769, 32'd7581},
{32'd8748, -32'd5884, 32'd9809, 32'd689},
{32'd591, 32'd8415, 32'd269, -32'd12594},
{-32'd10879, 32'd24977, -32'd4960, -32'd5571},
{-32'd5046, -32'd8548, -32'd2236, 32'd9024},
{32'd4530, 32'd6242, 32'd11425, -32'd630},
{32'd2697, 32'd7272, -32'd554, 32'd1827},
{32'd3171, 32'd33, 32'd9040, -32'd9985},
{32'd5861, 32'd18990, 32'd1479, 32'd3183},
{32'd3011, -32'd14656, -32'd3218, -32'd2518},
{-32'd8792, -32'd19014, -32'd70, 32'd1526},
{32'd955, 32'd5920, -32'd10028, -32'd5069},
{32'd4063, -32'd13882, 32'd843, 32'd6491},
{-32'd2198, 32'd2877, -32'd1486, -32'd3097},
{32'd1873, -32'd1385, -32'd12271, -32'd597},
{32'd2040, 32'd13468, -32'd282, 32'd7645},
{32'd7039, 32'd6774, 32'd6072, -32'd9293},
{32'd4802, 32'd3950, -32'd6877, 32'd736},
{-32'd13167, -32'd4201, -32'd1235, -32'd10926},
{32'd970, 32'd3403, 32'd45, 32'd2302},
{32'd7926, 32'd7140, 32'd8902, -32'd2796},
{32'd5101, 32'd1014, -32'd2493, 32'd4478},
{-32'd3606, -32'd10658, 32'd5613, 32'd4178},
{-32'd6212, -32'd3029, -32'd3133, -32'd5930},
{32'd382, -32'd13377, -32'd2824, 32'd14404},
{-32'd2577, -32'd12150, -32'd14187, -32'd4459},
{32'd566, -32'd9819, 32'd5481, 32'd8584},
{-32'd4230, -32'd9836, -32'd1638, 32'd1749},
{32'd4081, -32'd1716, 32'd9652, -32'd17751},
{32'd3692, -32'd1968, -32'd2752, 32'd9403},
{-32'd597, -32'd2786, 32'd6675, -32'd4282},
{32'd3715, -32'd13612, -32'd8355, -32'd1154},
{-32'd972, -32'd5842, -32'd19864, -32'd11165},
{-32'd4026, 32'd2812, 32'd6404, 32'd6686},
{32'd229, 32'd14729, 32'd4724, 32'd1367},
{-32'd3745, -32'd5054, -32'd3719, -32'd1281},
{-32'd4369, -32'd3311, -32'd7469, 32'd3196},
{32'd1213, -32'd265, 32'd7143, 32'd10584},
{-32'd3760, -32'd9329, -32'd3232, -32'd4640},
{-32'd1518, -32'd15123, -32'd19641, 32'd4341},
{32'd1084, -32'd13128, -32'd10212, -32'd4702},
{-32'd13948, -32'd7723, 32'd13371, 32'd12783},
{-32'd1556, 32'd7834, 32'd371, -32'd2216},
{-32'd14870, -32'd786, -32'd1488, 32'd15448},
{32'd6627, -32'd10669, -32'd15317, -32'd4233},
{32'd8838, 32'd3087, -32'd6725, -32'd8748},
{-32'd4732, 32'd1787, 32'd4629, -32'd7979},
{-32'd11053, 32'd3036, 32'd7035, 32'd7966},
{-32'd11221, -32'd13938, -32'd4513, -32'd16148},
{32'd6193, 32'd10564, 32'd11408, 32'd8962},
{32'd2675, 32'd14705, -32'd8759, -32'd3019},
{32'd11021, 32'd5265, 32'd5817, 32'd13267},
{-32'd13773, -32'd3815, -32'd1854, -32'd88},
{-32'd1097, 32'd12284, 32'd2232, -32'd8323},
{32'd15171, -32'd6429, 32'd5999, -32'd19900},
{-32'd6781, 32'd17590, 32'd6903, -32'd8316},
{-32'd7362, -32'd10917, -32'd5738, 32'd8811},
{32'd1860, -32'd5760, -32'd13998, 32'd20759},
{-32'd146, 32'd16080, 32'd4673, 32'd1006},
{-32'd10269, -32'd815, 32'd1575, -32'd2011},
{-32'd2742, -32'd7377, -32'd1592, 32'd11610},
{32'd202, -32'd4199, -32'd7528, -32'd3972},
{32'd2106, 32'd11776, 32'd7054, 32'd13211},
{-32'd535, -32'd6717, 32'd7268, 32'd12759},
{32'd2081, 32'd7516, 32'd443, -32'd7455},
{32'd10197, -32'd5933, -32'd6121, 32'd14899},
{32'd6410, -32'd9292, 32'd7157, 32'd10890},
{32'd7722, -32'd15614, -32'd2284, -32'd10078},
{-32'd8398, 32'd989, 32'd7233, 32'd3931},
{32'd7151, -32'd4917, -32'd3756, -32'd11361},
{-32'd4317, 32'd10195, -32'd8469, -32'd2566},
{32'd6358, -32'd2954, 32'd1886, 32'd648},
{-32'd4929, 32'd8961, 32'd5825, -32'd6939},
{-32'd2509, -32'd9737, -32'd2645, -32'd1013},
{-32'd784, -32'd10852, 32'd5045, 32'd5198},
{32'd3744, -32'd20408, -32'd5126, 32'd1654},
{-32'd4737, -32'd1899, 32'd6778, 32'd50},
{-32'd1095, -32'd6073, 32'd1323, -32'd5774},
{32'd1176, -32'd19903, 32'd8988, 32'd197},
{-32'd4650, 32'd962, -32'd5489, 32'd2253},
{32'd11290, -32'd758, -32'd859, 32'd3280},
{-32'd13050, -32'd12597, -32'd6459, 32'd5728},
{32'd6692, -32'd2288, -32'd9730, 32'd12225},
{32'd16473, 32'd12799, 32'd1588, -32'd9800},
{32'd7476, -32'd10020, -32'd12043, 32'd9467},
{-32'd1548, 32'd4012, 32'd9885, 32'd1494},
{32'd2330, -32'd6998, -32'd4884, 32'd2157},
{32'd696, -32'd4965, 32'd4136, 32'd18264},
{32'd3458, 32'd1644, -32'd11641, -32'd4293},
{-32'd8213, -32'd1453, 32'd10540, 32'd13256},
{-32'd5931, -32'd2298, -32'd463, -32'd14829},
{-32'd2556, 32'd8690, 32'd833, -32'd5437},
{32'd13193, -32'd10421, 32'd4261, 32'd223},
{-32'd5964, -32'd11801, -32'd5131, 32'd1261},
{-32'd3742, -32'd17811, 32'd3525, 32'd3662},
{-32'd2679, -32'd3759, -32'd994, 32'd895},
{-32'd838, -32'd3348, -32'd897, -32'd2467},
{32'd5042, -32'd4300, -32'd2199, 32'd2886},
{32'd496, -32'd3387, -32'd5585, -32'd3356},
{32'd6186, 32'd3167, 32'd5302, 32'd12219},
{-32'd3957, -32'd10476, -32'd18262, 32'd13144},
{-32'd11829, -32'd6534, 32'd7223, 32'd4393},
{-32'd2422, 32'd2632, 32'd2947, -32'd3256},
{32'd992, 32'd6974, 32'd3815, 32'd7452},
{-32'd155, 32'd1367, -32'd9632, 32'd2936},
{-32'd10352, 32'd6258, 32'd6564, -32'd6262},
{32'd1343, -32'd8967, -32'd7275, -32'd6082},
{32'd6980, 32'd9037, 32'd13699, 32'd7639},
{32'd8480, -32'd4467, -32'd633, -32'd694},
{-32'd6009, -32'd7761, 32'd8824, -32'd2168},
{-32'd4963, 32'd3774, 32'd7141, -32'd4641},
{-32'd5970, 32'd3103, 32'd8479, 32'd1514},
{-32'd2148, 32'd1044, -32'd3332, -32'd6664},
{32'd4995, -32'd12933, 32'd201, -32'd5975},
{-32'd1762, 32'd621, 32'd11413, 32'd8883},
{-32'd4994, 32'd13168, -32'd1284, -32'd3189},
{-32'd8206, -32'd6849, 32'd1244, 32'd6230},
{-32'd3140, -32'd7746, -32'd5511, 32'd173},
{32'd20920, -32'd4288, -32'd1363, 32'd14974},
{-32'd12172, -32'd7605, -32'd606, 32'd4011},
{-32'd13452, 32'd2327, -32'd736, 32'd139},
{-32'd1254, -32'd16868, -32'd11538, -32'd15380},
{-32'd3953, 32'd19525, -32'd5966, -32'd4515},
{32'd10337, 32'd8783, -32'd4629, 32'd3182},
{32'd4062, 32'd801, 32'd1751, 32'd17659},
{32'd9777, -32'd18638, -32'd12819, -32'd2907},
{32'd6325, 32'd6779, -32'd4424, -32'd10871},
{-32'd10583, -32'd8891, 32'd3385, -32'd5265},
{-32'd3555, -32'd435, -32'd2520, 32'd1667},
{-32'd4088, -32'd4226, -32'd18279, 32'd12104},
{32'd10156, 32'd751, 32'd2967, 32'd10940},
{-32'd7570, -32'd6090, 32'd5496, 32'd3383},
{-32'd7095, -32'd11972, -32'd8282, -32'd303},
{32'd10544, 32'd3732, -32'd14600, -32'd1368},
{-32'd6534, 32'd952, 32'd4883, -32'd754},
{32'd7398, -32'd9124, 32'd9933, -32'd12181},
{-32'd1176, -32'd18645, -32'd3343, 32'd7},
{-32'd2149, 32'd1304, 32'd12675, -32'd1300},
{32'd5471, -32'd2523, -32'd6559, -32'd543},
{32'd1950, 32'd2799, 32'd4841, -32'd1610},
{32'd6658, -32'd7828, 32'd5789, 32'd1467},
{-32'd12560, -32'd6819, 32'd13537, -32'd9126},
{-32'd3692, -32'd11543, -32'd16093, 32'd10700},
{-32'd13605, 32'd6672, 32'd1482, 32'd4594},
{-32'd1913, -32'd7595, 32'd12037, 32'd4165},
{32'd2553, -32'd2123, -32'd5150, -32'd980},
{-32'd6748, 32'd10121, -32'd24, -32'd405},
{32'd5280, -32'd3125, 32'd1102, -32'd12387},
{32'd749, -32'd3964, -32'd608, -32'd3696},
{32'd5611, 32'd2491, 32'd6800, 32'd837},
{-32'd5443, 32'd5475, 32'd17053, -32'd104},
{-32'd1358, 32'd6128, -32'd228, 32'd4936},
{-32'd1377, 32'd6215, 32'd9946, 32'd1306},
{-32'd1361, 32'd2721, 32'd16460, -32'd4873},
{-32'd3396, -32'd7719, -32'd1597, -32'd8356},
{-32'd3763, -32'd3892, 32'd900, -32'd21984},
{32'd1925, 32'd16400, 32'd1351, 32'd6947},
{-32'd2902, 32'd16549, -32'd2696, -32'd7863},
{-32'd2210, -32'd6965, 32'd4875, 32'd2527},
{32'd360, -32'd1202, -32'd2918, -32'd4633},
{32'd7567, 32'd2269, 32'd2229, -32'd2290},
{-32'd2241, 32'd904, 32'd9436, -32'd226},
{32'd6569, 32'd4230, 32'd4183, 32'd6979},
{-32'd8839, -32'd3427, -32'd12421, -32'd19937},
{-32'd3305, -32'd1609, -32'd4058, -32'd1870},
{-32'd573, 32'd15488, 32'd2888, 32'd2811},
{32'd941, 32'd6154, 32'd1049, 32'd23118},
{32'd19144, 32'd12128, -32'd26239, 32'd5617},
{32'd6982, 32'd7842, -32'd3309, -32'd6426},
{32'd10295, 32'd1247, 32'd4544, -32'd5206},
{32'd4029, 32'd11279, -32'd2509, -32'd9389},
{32'd723, -32'd2001, -32'd5439, 32'd367},
{32'd6277, 32'd6278, 32'd25, 32'd3662},
{-32'd5972, -32'd4956, 32'd6628, 32'd3708},
{32'd5967, -32'd13997, -32'd4901, -32'd11007},
{-32'd6511, 32'd6382, 32'd4131, 32'd7658},
{32'd1650, 32'd7001, 32'd11708, -32'd2428},
{32'd13440, 32'd3351, 32'd6168, 32'd14048},
{-32'd4143, -32'd8234, 32'd659, 32'd8173},
{32'd8462, 32'd3866, -32'd5887, -32'd14486},
{32'd5624, -32'd9245, -32'd4372, 32'd13453},
{-32'd929, -32'd3690, -32'd7368, 32'd8733},
{-32'd8033, -32'd15084, 32'd5483, 32'd2593},
{-32'd5538, 32'd6495, 32'd4223, 32'd4821},
{-32'd2585, 32'd17113, 32'd535, 32'd13269},
{32'd3826, -32'd10878, -32'd2357, -32'd10328}
},
{{32'd6378, 32'd10798, 32'd5019, 32'd11781},
{-32'd4771, -32'd4575, -32'd2961, 32'd2756},
{32'd7311, 32'd5790, 32'd11038, 32'd3955},
{-32'd6024, 32'd5797, -32'd1950, -32'd5217},
{32'd11575, 32'd2060, -32'd4194, -32'd6725},
{32'd3330, -32'd4558, -32'd5600, 32'd3131},
{32'd3562, 32'd2879, 32'd4267, 32'd2396},
{-32'd2597, -32'd8168, -32'd5361, -32'd8245},
{32'd4336, 32'd4911, 32'd5653, 32'd2938},
{32'd13296, 32'd6638, 32'd4383, 32'd7275},
{-32'd2088, -32'd6577, -32'd4137, 32'd430},
{32'd8896, 32'd5486, 32'd13468, 32'd3174},
{-32'd5444, -32'd5451, -32'd3841, 32'd6136},
{-32'd11204, -32'd6047, -32'd3983, -32'd11044},
{-32'd7970, 32'd1287, 32'd3655, -32'd9777},
{-32'd1916, -32'd8641, -32'd7302, -32'd2328},
{32'd5500, -32'd774, 32'd7521, -32'd2322},
{32'd5577, 32'd4842, 32'd11482, 32'd5921},
{32'd7922, -32'd596, -32'd2840, 32'd2496},
{32'd3721, -32'd1095, 32'd4282, -32'd8106},
{32'd9189, -32'd5425, -32'd560, 32'd445},
{-32'd12201, -32'd7828, -32'd2465, -32'd8399},
{-32'd1027, -32'd2560, -32'd5756, -32'd2334},
{-32'd239, -32'd1763, -32'd1463, 32'd832},
{32'd10929, 32'd1670, 32'd1233, 32'd4841},
{-32'd14188, -32'd731, -32'd6189, -32'd2124},
{32'd362, 32'd2086, 32'd3851, -32'd7234},
{-32'd9975, -32'd2605, 32'd4191, 32'd7351},
{32'd4235, -32'd8585, 32'd7345, 32'd2861},
{-32'd2170, 32'd2493, -32'd5244, 32'd7619},
{32'd1264, -32'd2169, 32'd4399, 32'd14791},
{-32'd18596, -32'd324, 32'd3621, -32'd2046},
{32'd8897, -32'd1969, -32'd690, 32'd719},
{-32'd8440, -32'd2020, -32'd3954, -32'd6716},
{32'd7261, 32'd5875, 32'd12118, 32'd4096},
{-32'd5403, -32'd4484, 32'd2756, -32'd2730},
{32'd864, -32'd6669, -32'd1621, -32'd2344},
{-32'd1209, -32'd266, 32'd2735, -32'd5797},
{32'd2995, 32'd11311, 32'd7908, -32'd1406},
{32'd1340, 32'd5392, 32'd8250, 32'd3132},
{32'd4057, 32'd8567, 32'd9959, -32'd1307},
{32'd10733, 32'd9115, -32'd432, 32'd9994},
{32'd5535, 32'd6260, 32'd23007, -32'd6354},
{-32'd4790, -32'd12438, -32'd3836, -32'd7731},
{-32'd4731, -32'd7967, -32'd10825, -32'd10222},
{32'd3051, -32'd9058, -32'd6628, -32'd403},
{32'd605, -32'd2704, -32'd11396, -32'd4865},
{-32'd2376, 32'd644, -32'd11576, -32'd17075},
{32'd7156, -32'd4056, -32'd1592, 32'd7015},
{32'd4360, -32'd6047, 32'd4913, -32'd5870},
{-32'd3708, 32'd1577, -32'd9583, -32'd7974},
{-32'd5305, 32'd5883, 32'd145, -32'd6023},
{-32'd3290, -32'd7152, -32'd352, 32'd2871},
{32'd1749, 32'd1610, -32'd3778, -32'd809},
{32'd12140, 32'd5314, 32'd4056, -32'd2567},
{-32'd1570, -32'd3972, -32'd4808, -32'd598},
{32'd5600, -32'd3631, -32'd5272, 32'd11702},
{-32'd2651, -32'd10186, -32'd18734, -32'd6429},
{-32'd5144, -32'd6174, -32'd3765, -32'd7093},
{32'd2086, -32'd1460, 32'd7130, -32'd3328},
{-32'd246, 32'd1366, 32'd4942, -32'd4635},
{-32'd8834, 32'd1423, 32'd3832, -32'd3323},
{-32'd6485, -32'd4068, -32'd5685, -32'd11169},
{-32'd1211, -32'd8356, -32'd2881, -32'd12343},
{-32'd5311, -32'd3184, 32'd2729, 32'd4556},
{32'd4519, 32'd5883, 32'd8026, 32'd5500},
{-32'd754, -32'd569, 32'd835, -32'd8929},
{-32'd11916, -32'd3342, -32'd748, -32'd4543},
{32'd8787, 32'd551, -32'd4036, 32'd2541},
{-32'd2178, 32'd98, 32'd6958, 32'd7140},
{-32'd8542, 32'd1543, -32'd7807, 32'd1496},
{-32'd1409, -32'd2812, 32'd5093, -32'd4062},
{-32'd1129, 32'd3967, -32'd4269, -32'd5055},
{-32'd430, -32'd5725, -32'd9365, 32'd1330},
{-32'd2266, 32'd6276, 32'd37, 32'd6406},
{32'd5820, -32'd1788, -32'd8377, -32'd8108},
{32'd4483, -32'd5452, -32'd1947, -32'd12405},
{32'd715, -32'd16487, -32'd4212, 32'd2094},
{32'd1653, 32'd6314, 32'd6829, 32'd8079},
{-32'd6837, -32'd3537, 32'd4543, -32'd4566},
{32'd7377, -32'd1098, 32'd4485, -32'd3556},
{32'd14732, -32'd10377, -32'd7366, 32'd9},
{32'd9345, -32'd11207, -32'd2432, -32'd10898},
{32'd2827, -32'd2711, 32'd16047, 32'd2249},
{-32'd4973, -32'd900, 32'd5229, -32'd11370},
{32'd136, -32'd787, -32'd4163, 32'd603},
{32'd5460, 32'd8728, 32'd5556, 32'd4146},
{-32'd5809, -32'd7278, -32'd10470, -32'd13396},
{-32'd5873, -32'd1746, 32'd9164, -32'd994},
{-32'd17381, 32'd1316, 32'd544, 32'd5809},
{32'd2161, 32'd4861, -32'd3416, 32'd8001},
{-32'd814, -32'd1009, 32'd2083, -32'd6536},
{-32'd4021, -32'd3358, -32'd3236, -32'd724},
{32'd3800, -32'd2386, 32'd2795, 32'd3309},
{-32'd8643, 32'd2268, 32'd3432, -32'd4386},
{-32'd2131, 32'd11570, 32'd5163, 32'd3563},
{32'd13869, 32'd4680, 32'd6686, -32'd2328},
{32'd6229, 32'd2453, 32'd1447, 32'd2748},
{32'd1528, -32'd1845, 32'd6333, 32'd6769},
{32'd1173, 32'd11400, 32'd8989, 32'd1329},
{-32'd4903, -32'd11878, 32'd2027, -32'd2935},
{32'd3390, -32'd6202, 32'd950, 32'd3346},
{32'd1113, 32'd3052, 32'd4070, -32'd4123},
{32'd4355, -32'd1562, 32'd625, 32'd3343},
{32'd10252, -32'd5409, 32'd3849, 32'd8580},
{-32'd9583, 32'd5182, 32'd3378, 32'd2829},
{32'd40, 32'd983, -32'd15459, 32'd12441},
{-32'd3627, -32'd5931, -32'd799, 32'd2649},
{32'd13725, -32'd881, 32'd8021, 32'd14649},
{-32'd5018, -32'd8130, -32'd998, -32'd4134},
{-32'd2977, -32'd8773, -32'd6510, -32'd12002},
{32'd10717, 32'd938, 32'd5232, -32'd7068},
{32'd5347, 32'd2936, 32'd763, -32'd3070},
{-32'd3386, 32'd3416, 32'd7687, -32'd431},
{32'd5256, 32'd1899, -32'd2933, -32'd3104},
{32'd3020, -32'd4025, 32'd8936, -32'd6298},
{32'd1604, -32'd592, -32'd3529, -32'd3404},
{-32'd9980, 32'd284, 32'd11551, -32'd4858},
{-32'd6022, -32'd7505, -32'd3238, -32'd5431},
{32'd10323, 32'd14472, 32'd4429, 32'd9199},
{-32'd10056, 32'd9910, 32'd2973, 32'd5673},
{-32'd343, 32'd1893, 32'd3861, -32'd4383},
{-32'd4984, 32'd1750, -32'd4451, -32'd5179},
{-32'd3007, 32'd3417, 32'd3957, 32'd7799},
{32'd2190, 32'd10072, 32'd11526, -32'd2591},
{-32'd1620, 32'd2892, -32'd5282, 32'd13282},
{32'd1529, -32'd192, -32'd15296, -32'd543},
{-32'd3275, -32'd5788, -32'd2238, -32'd14622},
{-32'd3492, 32'd4475, 32'd1164, 32'd13387},
{-32'd1575, -32'd11050, -32'd6379, 32'd141},
{-32'd7118, -32'd1173, -32'd214, -32'd1199},
{-32'd2436, -32'd2281, 32'd3329, -32'd9841},
{-32'd5215, -32'd16090, 32'd329, -32'd4903},
{-32'd4338, 32'd5503, 32'd3819, -32'd6418},
{32'd3266, 32'd814, -32'd4622, -32'd7790},
{32'd2303, -32'd16744, -32'd6153, 32'd1882},
{32'd4704, 32'd8077, -32'd10857, -32'd2501},
{-32'd641, 32'd9556, -32'd3404, 32'd9790},
{32'd1166, 32'd4722, 32'd18196, 32'd956},
{32'd2960, -32'd1773, -32'd4998, -32'd8207},
{32'd1199, -32'd1066, -32'd7016, -32'd7022},
{32'd2802, -32'd339, -32'd5089, -32'd1607},
{-32'd1012, 32'd3952, -32'd7477, 32'd8368},
{32'd7802, -32'd1422, 32'd7546, -32'd3505},
{32'd5273, 32'd5849, 32'd11174, 32'd2953},
{32'd2791, 32'd6949, 32'd7692, 32'd536},
{-32'd10017, -32'd3530, -32'd1416, -32'd5422},
{32'd3287, 32'd1509, 32'd4907, 32'd3161},
{32'd188, 32'd4856, 32'd2406, 32'd351},
{32'd2217, -32'd647, 32'd10761, -32'd8943},
{32'd3510, -32'd433, -32'd2187, -32'd2364},
{32'd10173, 32'd4283, 32'd1403, -32'd6588},
{32'd1385, -32'd11733, -32'd906, 32'd3913},
{32'd4797, -32'd4347, 32'd1203, -32'd9399},
{-32'd6542, -32'd7053, -32'd9840, -32'd4047},
{32'd2031, 32'd5843, -32'd208, -32'd533},
{32'd7611, 32'd3147, 32'd3402, 32'd1329},
{32'd1093, -32'd710, 32'd2131, -32'd5294},
{-32'd2237, -32'd2551, -32'd4117, -32'd531},
{32'd8571, -32'd2055, 32'd3244, -32'd4338},
{32'd931, -32'd6647, -32'd731, -32'd6431},
{-32'd11762, -32'd3509, 32'd233, -32'd10362},
{32'd10630, -32'd9219, -32'd2956, -32'd2418},
{32'd2840, -32'd7146, 32'd4223, 32'd12080},
{32'd2179, 32'd8701, 32'd3244, 32'd5146},
{-32'd3210, -32'd3330, 32'd255, -32'd869},
{-32'd11600, -32'd1765, 32'd1648, 32'd3981},
{-32'd1853, -32'd11686, 32'd4470, -32'd3105},
{32'd3678, -32'd3356, -32'd6966, -32'd1690},
{-32'd957, 32'd5140, -32'd3139, 32'd4556},
{-32'd8185, 32'd2895, 32'd1986, 32'd1287},
{-32'd5432, -32'd2306, -32'd7193, -32'd5832},
{32'd2004, 32'd7268, 32'd9107, 32'd8267},
{-32'd3826, 32'd79, -32'd5695, 32'd2012},
{32'd6970, 32'd2964, -32'd12235, 32'd6641},
{-32'd2663, -32'd11005, 32'd2337, 32'd1596},
{32'd29, 32'd9998, -32'd66, -32'd6221},
{32'd1845, 32'd1791, -32'd13760, 32'd7696},
{32'd444, -32'd4190, -32'd8286, -32'd3214},
{-32'd10016, -32'd1700, -32'd6037, -32'd8293},
{-32'd3057, -32'd6370, -32'd6740, -32'd3839},
{-32'd5554, -32'd10978, -32'd11372, -32'd6882},
{32'd4079, -32'd7903, -32'd8587, 32'd3634},
{-32'd869, -32'd5119, -32'd12232, 32'd1178},
{-32'd11169, -32'd9660, -32'd694, 32'd121},
{-32'd400, 32'd8159, 32'd4809, 32'd14983},
{-32'd2751, 32'd2152, 32'd4321, 32'd5324},
{-32'd488, 32'd2911, 32'd4460, 32'd1841},
{-32'd3679, -32'd6250, 32'd5103, -32'd2129},
{-32'd798, -32'd4412, -32'd10112, -32'd7234},
{32'd3012, 32'd1351, 32'd1794, 32'd702},
{-32'd7340, -32'd1907, -32'd11265, 32'd2847},
{-32'd2188, 32'd6465, -32'd6984, 32'd10891},
{-32'd973, 32'd5301, 32'd6156, 32'd8487},
{-32'd7029, 32'd4261, 32'd2225, 32'd9364},
{32'd1113, -32'd6602, 32'd5123, -32'd692},
{-32'd1444, 32'd2554, -32'd1170, 32'd1419},
{32'd4445, -32'd1155, 32'd5728, 32'd2407},
{32'd5634, 32'd11322, -32'd22067, 32'd1936},
{32'd9884, 32'd4049, 32'd1633, 32'd4309},
{-32'd5722, -32'd10003, -32'd14749, -32'd3359},
{-32'd3983, 32'd608, 32'd3991, -32'd4420},
{32'd297, -32'd1763, 32'd1521, 32'd1522},
{32'd4156, 32'd1814, 32'd11846, -32'd2870},
{-32'd6696, -32'd4310, -32'd3179, -32'd1414},
{32'd3570, 32'd8385, 32'd5120, 32'd2609},
{32'd6232, -32'd3704, -32'd7262, 32'd6796},
{-32'd2920, 32'd2552, -32'd2811, 32'd3137},
{32'd580, 32'd3270, -32'd2844, -32'd1406},
{32'd2637, 32'd5751, 32'd12992, -32'd1166},
{32'd9853, 32'd8194, -32'd13558, -32'd10601},
{32'd6019, 32'd6967, -32'd272, 32'd4935},
{-32'd11154, 32'd9296, -32'd298, -32'd7536},
{-32'd6579, -32'd7690, 32'd6715, 32'd4768},
{32'd3081, 32'd980, -32'd2205, -32'd9488},
{-32'd6911, -32'd2210, 32'd1201, -32'd4046},
{-32'd6270, 32'd5371, -32'd4140, -32'd1554},
{-32'd2360, 32'd2274, 32'd1149, -32'd2877},
{32'd671, 32'd9881, 32'd7502, 32'd3030},
{-32'd2759, 32'd3245, 32'd2615, -32'd2529},
{-32'd1065, -32'd730, -32'd5528, 32'd1808},
{-32'd3522, -32'd3924, 32'd1723, 32'd292},
{32'd20418, 32'd1141, 32'd521, -32'd405},
{32'd3969, -32'd761, -32'd3692, 32'd10082},
{32'd4161, 32'd673, 32'd913, 32'd1614},
{32'd1819, -32'd6634, 32'd5053, -32'd3755},
{-32'd6835, -32'd5282, -32'd3903, -32'd6951},
{-32'd6243, -32'd2450, 32'd36, -32'd435},
{32'd3421, 32'd9854, -32'd6533, -32'd1522},
{-32'd6868, 32'd5965, -32'd1331, -32'd530},
{-32'd9299, 32'd4793, 32'd8687, -32'd4698},
{-32'd8987, 32'd11226, 32'd11985, -32'd8440},
{-32'd582, 32'd5353, -32'd10281, 32'd2245},
{32'd4735, 32'd1442, -32'd849, -32'd10730},
{-32'd10044, -32'd6923, 32'd4283, -32'd13097},
{-32'd3385, -32'd1066, -32'd1693, -32'd13901},
{-32'd6175, 32'd3233, 32'd7560, -32'd1408},
{-32'd4727, -32'd3779, 32'd5358, -32'd1159},
{32'd8047, -32'd650, -32'd2410, -32'd886},
{-32'd10477, 32'd4499, -32'd46, 32'd3842},
{32'd2662, 32'd1947, -32'd2285, 32'd10150},
{32'd3685, 32'd8945, 32'd891, -32'd3606},
{-32'd10730, -32'd4869, -32'd2149, -32'd9151},
{-32'd6149, 32'd3970, -32'd11675, 32'd7429},
{32'd6538, 32'd2979, 32'd1547, 32'd1610},
{32'd5607, 32'd1705, 32'd8414, -32'd11337},
{-32'd8685, 32'd1750, 32'd3508, -32'd856},
{-32'd3752, 32'd272, 32'd1599, 32'd10738},
{-32'd2643, 32'd5219, -32'd1415, 32'd2552},
{-32'd9889, -32'd2041, 32'd12113, -32'd1091},
{32'd3479, -32'd5668, -32'd5005, -32'd1373},
{-32'd8536, -32'd3131, -32'd5437, 32'd294},
{-32'd414, -32'd1783, -32'd3144, 32'd656},
{-32'd909, -32'd2451, 32'd2178, -32'd1752},
{-32'd2266, -32'd4651, -32'd2722, -32'd10749},
{-32'd1918, 32'd8883, -32'd238, 32'd14153},
{-32'd3172, -32'd7252, -32'd6385, -32'd9414},
{-32'd5933, 32'd1299, 32'd3660, -32'd12391},
{-32'd5637, -32'd7479, -32'd5096, -32'd13848},
{32'd1617, 32'd4865, 32'd3617, 32'd3941},
{-32'd3533, -32'd3352, -32'd620, 32'd7247},
{32'd12409, 32'd2890, -32'd3840, 32'd3568},
{32'd2996, -32'd8752, -32'd2422, -32'd3027},
{-32'd4765, 32'd2071, -32'd4976, 32'd9251},
{-32'd7851, 32'd4963, 32'd829, -32'd972},
{-32'd1614, -32'd8177, -32'd11246, 32'd5081},
{32'd1722, -32'd932, -32'd5693, 32'd10797},
{32'd3588, 32'd9448, -32'd784, 32'd161},
{-32'd5503, -32'd6523, -32'd5639, 32'd2655},
{-32'd3551, -32'd10086, -32'd5305, 32'd5110},
{32'd6353, 32'd7726, -32'd1088, -32'd5132},
{32'd6692, 32'd11947, 32'd4524, 32'd164},
{-32'd1489, -32'd10102, -32'd716, -32'd210},
{-32'd4109, -32'd4667, 32'd1078, -32'd6140},
{-32'd938, -32'd1244, 32'd4103, -32'd9259},
{-32'd3209, -32'd13226, 32'd2176, -32'd9708},
{32'd13666, 32'd7172, 32'd6428, 32'd8091},
{32'd308, 32'd962, -32'd3652, 32'd11281},
{-32'd2096, -32'd7979, 32'd220, -32'd8636},
{-32'd4580, -32'd2201, 32'd5494, 32'd9263},
{32'd7316, 32'd5997, 32'd8387, -32'd1879},
{-32'd941, -32'd1168, 32'd8888, 32'd6223},
{32'd4858, 32'd9336, 32'd4713, 32'd6597},
{-32'd3703, 32'd1320, -32'd5800, 32'd9589},
{32'd14124, 32'd9775, 32'd1545, 32'd1146},
{-32'd12250, -32'd4007, -32'd5725, -32'd11325},
{-32'd2411, 32'd1596, 32'd1874, 32'd5574},
{-32'd7190, -32'd3762, -32'd294, -32'd2148},
{32'd5969, -32'd3236, 32'd7162, -32'd4210},
{32'd2941, 32'd4268, 32'd1065, -32'd7602},
{32'd561, -32'd6260, -32'd9329, 32'd1843},
{32'd4250, 32'd4015, 32'd2590, 32'd5167},
{-32'd6015, -32'd1480, -32'd6828, -32'd4522},
{-32'd1406, 32'd3108, -32'd6209, 32'd1298},
{-32'd4960, 32'd3842, -32'd7569, -32'd184},
{32'd987, 32'd5256, -32'd7874, -32'd610},
{-32'd930, 32'd3566, -32'd3631, -32'd4413},
{32'd6275, 32'd3560, 32'd7504, -32'd4734},
{32'd6853, 32'd9304, 32'd2664, 32'd10786},
{-32'd5198, -32'd8440, 32'd1162, -32'd3558}
},
{{-32'd763, -32'd11635, -32'd7035, -32'd305},
{32'd1312, 32'd1021, -32'd10565, -32'd1675},
{-32'd9608, 32'd1474, 32'd5108, -32'd6761},
{-32'd1795, -32'd4869, 32'd676, 32'd10669},
{32'd678, -32'd3474, -32'd6797, 32'd5763},
{-32'd15650, -32'd8391, -32'd5165, 32'd1597},
{32'd8153, 32'd9836, -32'd791, -32'd4820},
{32'd3450, -32'd966, 32'd8139, 32'd3906},
{-32'd5563, 32'd9790, -32'd9379, 32'd10556},
{32'd9886, 32'd4657, 32'd3448, 32'd303},
{-32'd8081, 32'd3283, -32'd11929, 32'd2538},
{32'd605, -32'd353, -32'd1316, 32'd6036},
{-32'd6007, -32'd6034, -32'd10670, -32'd4358},
{-32'd1033, -32'd9359, 32'd6116, -32'd2104},
{-32'd14895, -32'd5645, 32'd8134, 32'd5},
{-32'd457, -32'd3742, -32'd11284, -32'd2416},
{32'd9402, -32'd3589, -32'd2635, -32'd5219},
{32'd16685, -32'd5830, -32'd2873, 32'd3987},
{32'd8160, -32'd14011, 32'd2173, 32'd11638},
{32'd11434, -32'd12177, 32'd10592, 32'd9668},
{-32'd981, 32'd12765, 32'd2170, 32'd3652},
{-32'd4881, -32'd10763, -32'd3246, 32'd5968},
{32'd9194, -32'd4311, 32'd6359, -32'd2854},
{-32'd1935, -32'd3342, 32'd3236, 32'd607},
{32'd5926, -32'd224, 32'd1329, -32'd7627},
{32'd2289, -32'd14436, 32'd1779, 32'd14020},
{32'd6758, -32'd11095, -32'd5711, -32'd2054},
{32'd9073, 32'd14456, 32'd9755, 32'd1891},
{32'd2035, 32'd3310, 32'd4750, 32'd889},
{32'd1932, 32'd3293, -32'd7832, 32'd4851},
{32'd6431, -32'd8685, 32'd12559, -32'd2302},
{-32'd15120, -32'd8480, 32'd8853, 32'd6478},
{32'd12778, -32'd11407, -32'd4298, -32'd1754},
{32'd12688, -32'd10187, -32'd7905, -32'd5104},
{32'd7322, 32'd11231, -32'd974, -32'd6530},
{-32'd3489, 32'd7730, -32'd9329, 32'd17},
{32'd3842, -32'd11054, 32'd6923, 32'd3565},
{32'd2128, 32'd10627, -32'd5412, -32'd86},
{32'd18045, -32'd1237, 32'd6942, -32'd2962},
{32'd5428, -32'd14450, -32'd5078, -32'd5449},
{-32'd8732, 32'd1890, 32'd9960, -32'd300},
{32'd8108, 32'd947, -32'd24645, -32'd1319},
{32'd9645, 32'd2535, 32'd7341, 32'd3782},
{32'd1594, -32'd6647, -32'd4042, -32'd5137},
{-32'd6178, 32'd4649, 32'd1257, -32'd6753},
{-32'd2887, 32'd12365, -32'd4788, -32'd475},
{-32'd7300, 32'd9177, -32'd1509, 32'd3346},
{-32'd6547, -32'd6814, -32'd4828, -32'd5245},
{32'd21558, -32'd2053, -32'd4489, -32'd6719},
{32'd1066, -32'd14747, -32'd10255, 32'd6892},
{-32'd4393, 32'd921, -32'd10086, -32'd4621},
{32'd3833, -32'd6800, -32'd746, -32'd2555},
{-32'd12798, -32'd5098, -32'd4074, -32'd3402},
{32'd15475, -32'd5885, 32'd7925, 32'd4682},
{32'd8541, -32'd4180, -32'd5593, 32'd6579},
{-32'd4547, -32'd1090, 32'd9665, -32'd4063},
{32'd9428, -32'd1062, -32'd11468, 32'd4538},
{32'd1843, -32'd5351, -32'd2558, -32'd7605},
{32'd2571, -32'd4043, 32'd7699, -32'd3553},
{32'd1141, -32'd4319, -32'd5806, -32'd7324},
{32'd2065, -32'd1896, 32'd8086, 32'd13281},
{-32'd12718, 32'd3658, 32'd11586, 32'd945},
{32'd3711, -32'd1268, 32'd3612, 32'd2956},
{-32'd1386, 32'd5822, 32'd3700, 32'd4660},
{32'd7439, -32'd4793, 32'd10885, -32'd8316},
{32'd9739, 32'd4379, -32'd6524, -32'd2426},
{32'd2083, -32'd3999, 32'd6017, 32'd2360},
{-32'd5895, -32'd3075, 32'd467, 32'd158},
{32'd7229, -32'd11292, -32'd1686, 32'd7071},
{32'd4215, 32'd13606, 32'd2339, -32'd3268},
{-32'd14212, -32'd2503, -32'd11197, 32'd3802},
{-32'd5902, 32'd2742, -32'd15758, -32'd7873},
{-32'd18, -32'd2662, -32'd11130, -32'd2130},
{-32'd1602, -32'd1713, 32'd248, 32'd9466},
{-32'd1684, 32'd8684, 32'd2209, 32'd6673},
{32'd3, 32'd1889, -32'd3361, -32'd1647},
{-32'd2106, -32'd3810, -32'd505, 32'd3147},
{-32'd1589, -32'd6265, -32'd6149, 32'd1366},
{32'd13443, 32'd5005, -32'd2279, -32'd589},
{-32'd10241, -32'd430, -32'd7191, -32'd8950},
{32'd3880, -32'd5859, 32'd4878, 32'd9306},
{32'd7615, -32'd6286, -32'd1324, -32'd2156},
{-32'd4273, 32'd183, 32'd2715, 32'd8948},
{32'd2774, -32'd6798, -32'd11043, 32'd2640},
{-32'd4181, -32'd14148, -32'd2502, 32'd5880},
{32'd10313, 32'd9308, 32'd13032, -32'd4500},
{32'd6281, -32'd13375, 32'd12573, 32'd3584},
{32'd2835, -32'd5031, -32'd2876, 32'd4154},
{-32'd9466, -32'd4091, -32'd277, -32'd3233},
{32'd3285, 32'd2399, 32'd6805, -32'd3874},
{32'd7369, -32'd15908, 32'd4442, -32'd2459},
{-32'd5938, 32'd11670, -32'd16273, 32'd13806},
{32'd2922, -32'd2297, 32'd1322, 32'd6421},
{-32'd2481, -32'd93, 32'd7466, 32'd6740},
{-32'd3187, 32'd6048, 32'd6208, 32'd914},
{-32'd6962, -32'd1204, -32'd2394, 32'd9785},
{32'd3505, -32'd6285, 32'd4295, 32'd7722},
{-32'd8788, 32'd4145, -32'd4008, -32'd1783},
{-32'd1301, 32'd52, 32'd2630, -32'd4260},
{32'd1357, 32'd6711, -32'd5123, -32'd2149},
{-32'd12056, 32'd2121, 32'd1024, 32'd4306},
{32'd11784, 32'd1901, -32'd2203, 32'd104},
{-32'd3183, 32'd1639, 32'd15730, 32'd4184},
{32'd594, 32'd13485, -32'd6624, -32'd1474},
{32'd5115, 32'd5437, 32'd1322, -32'd7168},
{-32'd7215, -32'd4924, -32'd3319, 32'd4890},
{-32'd8057, -32'd4518, 32'd1412, -32'd3230},
{32'd12871, 32'd9107, 32'd12820, 32'd8931},
{32'd5719, 32'd3893, 32'd1940, -32'd3357},
{32'd1659, 32'd2600, -32'd9457, -32'd3377},
{32'd6153, 32'd11467, -32'd4279, -32'd4935},
{32'd4342, 32'd1863, -32'd3983, -32'd8368},
{32'd8124, 32'd2158, -32'd14787, -32'd5334},
{32'd9207, -32'd3806, 32'd3485, 32'd4255},
{-32'd7632, -32'd7415, -32'd7670, 32'd3682},
{32'd1787, -32'd3202, 32'd2473, -32'd1003},
{32'd5514, 32'd4672, 32'd1977, -32'd5067},
{32'd12794, 32'd572, -32'd4897, 32'd6088},
{32'd3793, 32'd13010, 32'd8781, -32'd6757},
{32'd1758, 32'd13251, -32'd8787, 32'd1079},
{32'd4902, 32'd5286, 32'd3552, 32'd510},
{32'd4250, 32'd4209, 32'd2412, 32'd5237},
{32'd6333, 32'd5893, -32'd12781, -32'd10375},
{-32'd2976, 32'd558, 32'd5319, -32'd1174},
{-32'd11046, -32'd13190, -32'd7552, 32'd2816},
{-32'd15380, 32'd8570, 32'd3803, 32'd10397},
{32'd4798, -32'd7251, -32'd4546, -32'd2202},
{-32'd4884, 32'd8084, 32'd10149, -32'd1102},
{-32'd5209, -32'd7659, -32'd291, 32'd154},
{32'd2025, -32'd7900, 32'd3575, -32'd8662},
{-32'd7549, 32'd973, 32'd7049, 32'd4024},
{32'd4987, -32'd14609, -32'd195, -32'd3469},
{-32'd15173, -32'd3261, 32'd4022, 32'd4011},
{-32'd3771, 32'd4273, -32'd9674, 32'd5083},
{-32'd2278, 32'd6605, 32'd5368, 32'd5688},
{32'd8622, -32'd753, -32'd10654, -32'd7288},
{-32'd3577, 32'd249, -32'd8580, 32'd141},
{32'd3910, 32'd3339, -32'd10340, -32'd2655},
{32'd19452, 32'd15827, 32'd16484, 32'd4741},
{32'd528, -32'd122, 32'd11091, 32'd3306},
{-32'd6474, 32'd914, 32'd3688, 32'd4766},
{32'd2682, 32'd3065, 32'd692, 32'd765},
{-32'd8388, -32'd3092, 32'd2604, 32'd4750},
{-32'd12700, -32'd8367, 32'd2835, 32'd11872},
{32'd6031, -32'd3570, 32'd5429, 32'd700},
{32'd974, 32'd309, 32'd12022, 32'd2885},
{32'd544, -32'd11857, 32'd1084, 32'd10980},
{-32'd784, -32'd3429, -32'd6592, -32'd2850},
{-32'd7516, 32'd13718, 32'd7119, 32'd11645},
{-32'd14797, -32'd1192, -32'd2852, 32'd4833},
{32'd606, -32'd9013, 32'd1311, -32'd1157},
{32'd3043, -32'd2903, 32'd12196, 32'd6850},
{32'd4885, -32'd2693, -32'd9944, -32'd4007},
{-32'd7421, 32'd6701, -32'd2551, 32'd3713},
{-32'd3096, 32'd2672, -32'd2824, 32'd5273},
{-32'd8459, -32'd12266, 32'd7650, -32'd6466},
{32'd8682, -32'd6973, -32'd6608, 32'd5341},
{32'd1924, -32'd1710, 32'd11755, 32'd5923},
{-32'd7635, -32'd1288, 32'd5683, -32'd4206},
{32'd5448, -32'd3088, -32'd4332, 32'd9679},
{-32'd7376, 32'd2075, 32'd9423, 32'd11210},
{-32'd1462, -32'd4459, 32'd8939, -32'd5996},
{32'd3365, -32'd6537, 32'd6280, -32'd5811},
{32'd596, 32'd6719, 32'd12168, 32'd6591},
{-32'd5779, 32'd1210, -32'd9880, 32'd5138},
{-32'd5037, -32'd3402, -32'd4269, -32'd3890},
{-32'd11201, 32'd2728, 32'd3490, -32'd180},
{32'd7241, -32'd8267, -32'd3574, -32'd5132},
{32'd2608, -32'd7312, -32'd18276, -32'd2941},
{-32'd1263, -32'd3559, 32'd9537, 32'd1005},
{-32'd6632, 32'd5234, 32'd9113, 32'd5134},
{32'd13008, 32'd8640, -32'd3527, 32'd432},
{32'd13695, 32'd9899, -32'd7669, -32'd9318},
{32'd6406, 32'd9052, 32'd936, 32'd8391},
{32'd2810, 32'd2418, -32'd43, 32'd379},
{32'd3191, -32'd12301, -32'd4723, -32'd1255},
{-32'd2130, 32'd1694, 32'd10137, 32'd5287},
{-32'd4623, -32'd928, -32'd7673, -32'd6411},
{-32'd10802, -32'd2846, -32'd1389, 32'd333},
{-32'd8775, -32'd2029, -32'd3340, -32'd5480},
{-32'd2624, 32'd7269, 32'd8727, 32'd3510},
{-32'd5772, -32'd9033, 32'd108, -32'd1133},
{32'd866, -32'd7721, -32'd18728, -32'd9022},
{-32'd7660, -32'd3047, -32'd5779, -32'd646},
{32'd3609, -32'd13439, 32'd6926, 32'd3328},
{32'd83, 32'd2180, 32'd8513, -32'd10029},
{32'd2656, 32'd7452, 32'd561, 32'd776},
{-32'd5267, 32'd7465, -32'd10309, -32'd9811},
{-32'd496, 32'd7704, 32'd3771, 32'd8967},
{32'd3479, -32'd3827, 32'd1092, -32'd13379},
{-32'd6638, -32'd4474, 32'd1359, -32'd3292},
{-32'd6405, -32'd4312, -32'd15378, -32'd4431},
{32'd1583, 32'd220, 32'd444, -32'd2195},
{-32'd298, -32'd1899, 32'd5070, -32'd740},
{32'd5040, 32'd23739, -32'd3886, -32'd367},
{32'd13682, -32'd3513, 32'd1775, -32'd10710},
{-32'd3242, 32'd4889, -32'd5747, -32'd2768},
{32'd6359, -32'd2919, -32'd6687, -32'd2213},
{32'd4845, 32'd9187, 32'd5174, -32'd5840},
{32'd9963, -32'd1758, -32'd5608, -32'd1957},
{-32'd7297, -32'd9436, 32'd5592, -32'd3115},
{-32'd585, 32'd8942, 32'd3730, 32'd3747},
{-32'd2320, -32'd7032, -32'd2751, 32'd3704},
{32'd6671, -32'd2281, 32'd6728, -32'd1584},
{32'd5435, -32'd11819, 32'd4164, 32'd15617},
{32'd4372, 32'd5565, 32'd4794, -32'd2421},
{32'd10701, 32'd9057, -32'd712, 32'd2529},
{-32'd10755, -32'd1728, 32'd5371, 32'd4738},
{-32'd4293, 32'd2909, 32'd2765, -32'd1984},
{-32'd1647, 32'd6577, -32'd8017, 32'd303},
{-32'd3321, 32'd9029, -32'd15273, -32'd965},
{32'd12809, -32'd175, -32'd2847, -32'd7002},
{32'd8169, 32'd420, -32'd1038, 32'd1132},
{32'd685, 32'd13377, 32'd919, 32'd1036},
{-32'd8721, -32'd12491, -32'd6607, 32'd3871},
{-32'd5898, -32'd18795, 32'd4165, -32'd6020},
{32'd6673, 32'd12139, 32'd9160, 32'd25},
{32'd3009, 32'd4214, -32'd656, 32'd5581},
{-32'd2810, 32'd2551, 32'd12280, -32'd6177},
{-32'd2509, 32'd6802, -32'd528, -32'd10951},
{32'd891, 32'd4947, -32'd8788, -32'd3328},
{32'd3743, 32'd15104, 32'd2373, -32'd2074},
{32'd6907, 32'd3605, -32'd3836, 32'd3477},
{32'd482, -32'd2793, 32'd1619, -32'd2753},
{-32'd3338, -32'd15403, -32'd11389, -32'd939},
{32'd3238, 32'd2630, 32'd1384, 32'd5448},
{32'd11926, -32'd8096, 32'd11257, 32'd3834},
{-32'd7693, -32'd4611, -32'd2939, -32'd5067},
{32'd1958, -32'd4806, 32'd4762, -32'd134},
{32'd2328, 32'd4005, -32'd15334, -32'd5531},
{-32'd6929, 32'd381, -32'd12498, 32'd5446},
{-32'd2879, -32'd3699, 32'd140, 32'd413},
{-32'd6223, 32'd14894, -32'd8179, 32'd2264},
{-32'd6241, 32'd9183, -32'd7951, -32'd6060},
{32'd4577, -32'd9927, 32'd3345, -32'd4926},
{32'd1365, 32'd3533, 32'd7791, -32'd7847},
{-32'd3543, 32'd698, 32'd8020, 32'd5151},
{-32'd9536, -32'd1054, -32'd2741, -32'd7241},
{32'd3430, 32'd11862, -32'd11503, -32'd6118},
{-32'd11282, 32'd13317, -32'd3450, 32'd6747},
{32'd3024, 32'd2151, -32'd6260, -32'd3310},
{-32'd10191, 32'd4776, -32'd5357, 32'd9869},
{-32'd4388, 32'd12, 32'd9162, 32'd5351},
{-32'd5412, -32'd1615, -32'd12290, 32'd262},
{32'd5972, 32'd8725, -32'd6695, 32'd5298},
{-32'd7689, -32'd7372, 32'd4953, -32'd1396},
{-32'd4330, 32'd4118, -32'd5592, -32'd2840},
{-32'd3058, 32'd7519, 32'd4564, 32'd10836},
{-32'd810, 32'd4393, -32'd11055, -32'd468},
{-32'd321, 32'd9443, 32'd15009, 32'd29},
{32'd4153, -32'd6387, -32'd7156, -32'd3722},
{-32'd150, -32'd7803, 32'd8011, -32'd1277},
{32'd6349, -32'd12064, 32'd18529, -32'd854},
{-32'd14101, -32'd6858, 32'd12671, 32'd9176},
{32'd5008, -32'd3234, 32'd11120, 32'd7861},
{-32'd2010, 32'd2498, 32'd8222, 32'd2932},
{-32'd7031, -32'd1677, 32'd12601, 32'd10341},
{-32'd16844, -32'd530, 32'd2388, 32'd6315},
{32'd160, -32'd9742, -32'd1882, -32'd2514},
{32'd10986, 32'd9630, -32'd2018, -32'd4855},
{32'd4161, 32'd8424, 32'd14283, -32'd2717},
{-32'd5127, -32'd7859, 32'd2683, -32'd3652},
{-32'd10626, 32'd8180, 32'd272, -32'd5375},
{-32'd12091, -32'd3193, -32'd17675, -32'd5588},
{-32'd5568, 32'd9911, 32'd11792, 32'd4481},
{-32'd3448, 32'd12147, 32'd1812, 32'd9164},
{-32'd4404, -32'd6930, -32'd10626, -32'd9611},
{32'd8709, -32'd7695, -32'd11425, 32'd6048},
{32'd1804, 32'd3055, -32'd1752, 32'd1474},
{-32'd9442, 32'd11990, 32'd2487, 32'd571},
{-32'd3120, 32'd18068, -32'd3683, -32'd3302},
{32'd3981, 32'd3886, -32'd3704, -32'd3326},
{32'd2727, -32'd8794, 32'd6598, -32'd614},
{-32'd10990, 32'd18237, -32'd2053, -32'd3502},
{32'd2237, 32'd3767, -32'd2387, 32'd13864},
{32'd5223, -32'd66, -32'd6043, 32'd5683},
{32'd13224, 32'd8903, -32'd3317, -32'd140},
{-32'd2614, 32'd554, 32'd1267, 32'd4684},
{32'd1047, -32'd7332, 32'd803, -32'd3237},
{32'd11954, -32'd12744, 32'd1251, 32'd1630},
{32'd12243, 32'd11344, 32'd17536, 32'd3690},
{32'd2680, 32'd9092, -32'd2078, 32'd4451},
{-32'd1717, 32'd11006, 32'd5552, 32'd1774},
{-32'd1146, 32'd12481, -32'd16382, 32'd5251},
{32'd17296, 32'd2939, 32'd1216, 32'd1560},
{32'd866, -32'd10390, 32'd1511, -32'd3168},
{32'd10700, 32'd2046, 32'd4132, -32'd6139},
{32'd5355, 32'd75, 32'd3390, 32'd3387},
{32'd6613, 32'd13989, 32'd8270, -32'd4081},
{-32'd8116, 32'd8279, 32'd1934, -32'd13478},
{-32'd5659, -32'd3255, -32'd2677, 32'd760},
{-32'd10844, 32'd1716, -32'd5573, 32'd4403},
{-32'd1393, 32'd13349, 32'd1201, -32'd5441},
{-32'd3042, -32'd4236, -32'd11983, -32'd2204},
{-32'd1456, 32'd14959, -32'd4329, -32'd1623},
{32'd734, -32'd9406, -32'd11634, -32'd1985},
{-32'd5897, -32'd4180, 32'd5312, -32'd9344},
{32'd12923, -32'd5249, 32'd1031, 32'd1205},
{32'd2208, -32'd2130, 32'd133, 32'd1115},
{32'd1130, -32'd16357, -32'd6293, 32'd9063}
},
{{32'd1101, 32'd11698, 32'd7724, 32'd3826},
{32'd1981, 32'd1505, -32'd9530, 32'd145},
{32'd2881, 32'd1160, 32'd2648, 32'd1667},
{32'd2190, -32'd6931, -32'd1618, -32'd477},
{-32'd509, -32'd4409, 32'd1884, 32'd3744},
{-32'd12947, -32'd6950, 32'd6565, 32'd200},
{32'd5854, 32'd1640, -32'd8990, -32'd801},
{-32'd9823, 32'd2265, 32'd7960, 32'd1432},
{-32'd10790, -32'd5084, 32'd10213, -32'd9387},
{32'd2938, 32'd4941, 32'd615, 32'd5991},
{32'd8502, -32'd5275, 32'd3319, -32'd4440},
{-32'd197, 32'd9116, -32'd6306, -32'd3124},
{32'd1266, -32'd674, 32'd6003, 32'd7713},
{-32'd3830, -32'd1546, -32'd6125, -32'd494},
{-32'd2374, -32'd3019, -32'd14151, -32'd5057},
{32'd7976, -32'd403, -32'd4383, 32'd2858},
{32'd6656, 32'd4322, 32'd10302, 32'd7666},
{-32'd3196, 32'd1272, 32'd825, 32'd8763},
{-32'd590, -32'd2004, -32'd6182, -32'd509},
{32'd12359, 32'd2442, -32'd13343, -32'd5427},
{32'd2536, 32'd6675, -32'd6541, -32'd4616},
{32'd3600, 32'd3169, -32'd3693, -32'd1430},
{32'd188, -32'd381, -32'd1616, 32'd815},
{32'd2517, -32'd13032, -32'd2746, -32'd16467},
{32'd3674, 32'd11509, -32'd932, 32'd6577},
{32'd4165, -32'd8331, -32'd1959, -32'd3361},
{-32'd6741, 32'd1323, -32'd4790, -32'd5817},
{32'd7424, -32'd252, 32'd1454, -32'd1673},
{32'd15511, 32'd4344, 32'd3839, 32'd6122},
{-32'd1485, -32'd8765, 32'd6315, 32'd969},
{32'd8715, -32'd3449, -32'd1654, -32'd1544},
{-32'd4544, 32'd1389, -32'd2426, 32'd7293},
{-32'd1443, -32'd1051, 32'd4876, 32'd2187},
{-32'd6862, -32'd10261, -32'd8236, 32'd1228},
{32'd7888, 32'd10167, 32'd1462, 32'd8246},
{-32'd9168, -32'd5654, -32'd3653, -32'd1310},
{-32'd552, 32'd6526, 32'd6465, 32'd5648},
{32'd1688, 32'd2969, -32'd1995, -32'd3783},
{32'd11368, -32'd15242, -32'd3575, -32'd4219},
{-32'd14562, -32'd9140, -32'd5085, -32'd6031},
{-32'd175, 32'd14535, 32'd1358, 32'd3499},
{-32'd3116, -32'd514, -32'd2008, 32'd7750},
{32'd11229, 32'd706, -32'd1320, 32'd13040},
{-32'd514, 32'd1108, -32'd8012, 32'd4156},
{-32'd2992, 32'd3176, -32'd3509, -32'd8114},
{32'd11038, -32'd11095, -32'd7792, -32'd5958},
{-32'd2917, -32'd4577, -32'd7500, 32'd7640},
{-32'd6053, -32'd10924, -32'd3190, -32'd3115},
{32'd3751, 32'd3525, 32'd1222, -32'd8363},
{-32'd773, -32'd3388, -32'd7684, 32'd7713},
{-32'd1694, 32'd487, -32'd2270, -32'd135},
{-32'd9963, 32'd5091, 32'd2554, 32'd919},
{32'd3755, -32'd2389, 32'd5682, 32'd7079},
{-32'd6526, 32'd3793, -32'd870, 32'd3221},
{32'd12447, 32'd7901, -32'd9648, 32'd12680},
{32'd5334, 32'd3847, 32'd4688, -32'd1723},
{32'd3288, -32'd9423, 32'd2313, -32'd5958},
{-32'd4281, -32'd16324, -32'd5656, -32'd3131},
{32'd8739, -32'd2498, 32'd637, -32'd352},
{32'd6593, -32'd11387, -32'd5511, -32'd4292},
{-32'd10346, -32'd278, -32'd2195, -32'd8112},
{32'd5133, 32'd13746, 32'd1466, -32'd2876},
{-32'd3847, -32'd8388, -32'd2662, -32'd2095},
{32'd9206, -32'd2940, -32'd13286, 32'd7779},
{32'd1368, -32'd6845, -32'd3251, 32'd6249},
{32'd855, 32'd667, 32'd3315, 32'd7949},
{-32'd6317, 32'd1150, -32'd8064, -32'd2160},
{-32'd6762, -32'd7105, 32'd4564, -32'd12706},
{-32'd6749, 32'd178, -32'd9594, 32'd2418},
{-32'd1855, 32'd5188, 32'd5851, -32'd1065},
{-32'd7365, 32'd3640, -32'd1817, 32'd925},
{-32'd2233, -32'd8298, 32'd5619, 32'd8090},
{-32'd7748, -32'd4954, -32'd5087, 32'd4089},
{32'd10844, 32'd3662, -32'd5788, -32'd1526},
{32'd14602, 32'd3262, 32'd4522, 32'd717},
{-32'd2829, -32'd3690, -32'd2866, -32'd5425},
{32'd9847, -32'd2489, -32'd8670, -32'd1103},
{32'd6281, -32'd8801, -32'd6356, -32'd6671},
{32'd665, -32'd9641, 32'd6651, 32'd4964},
{-32'd5603, 32'd10126, -32'd678, 32'd4592},
{-32'd6103, 32'd4582, -32'd2951, -32'd6529},
{32'd4784, -32'd2976, 32'd1080, 32'd3885},
{32'd553, -32'd2481, 32'd1437, -32'd126},
{-32'd2520, 32'd8998, 32'd6872, 32'd8449},
{-32'd6656, -32'd6528, -32'd7488, 32'd7562},
{-32'd1821, -32'd5125, -32'd630, -32'd1156},
{32'd2094, -32'd1581, -32'd728, 32'd3579},
{32'd1385, -32'd6796, -32'd7075, -32'd6304},
{32'd750, -32'd3711, -32'd4484, -32'd8144},
{-32'd1978, -32'd9211, -32'd2652, 32'd839},
{32'd1684, -32'd3202, 32'd1544, 32'd10043},
{32'd1287, 32'd1452, -32'd9094, -32'd4973},
{-32'd5377, -32'd4851, -32'd4227, -32'd10240},
{32'd15124, 32'd10427, -32'd392, 32'd3467},
{32'd10948, -32'd1205, 32'd5449, 32'd6768},
{-32'd8467, 32'd6582, -32'd4193, 32'd8863},
{-32'd545, 32'd2937, -32'd203, 32'd4714},
{-32'd7753, 32'd9362, 32'd4202, 32'd6885},
{32'd7525, 32'd7593, 32'd3634, -32'd1530},
{-32'd1868, 32'd1916, 32'd2211, 32'd6793},
{-32'd688, -32'd6302, 32'd1782, 32'd1067},
{-32'd5688, -32'd2293, 32'd540, 32'd6843},
{-32'd321, 32'd3992, 32'd2868, 32'd2940},
{32'd8539, 32'd6878, 32'd9698, -32'd5098},
{32'd2596, 32'd393, 32'd953, 32'd9690},
{32'd7450, -32'd772, -32'd2772, -32'd2084},
{32'd3197, 32'd3766, 32'd11410, -32'd4135},
{-32'd3714, 32'd8863, 32'd915, -32'd2755},
{32'd10078, 32'd5376, -32'd11206, 32'd2431},
{32'd3841, -32'd3524, -32'd373, 32'd419},
{32'd2328, -32'd326, 32'd1885, -32'd2625},
{32'd4584, 32'd63, -32'd83, 32'd3731},
{32'd12338, 32'd4169, 32'd2668, 32'd1365},
{32'd106, 32'd10810, -32'd1814, -32'd9319},
{32'd8106, 32'd332, -32'd6688, 32'd8452},
{32'd1226, 32'd4950, -32'd4621, 32'd532},
{32'd13450, 32'd3430, 32'd6691, 32'd2912},
{-32'd5803, 32'd5502, 32'd2734, -32'd6584},
{-32'd18319, 32'd10357, -32'd1471, -32'd7853},
{32'd2674, 32'd2252, -32'd157, 32'd2356},
{-32'd209, 32'd6160, -32'd8948, 32'd4054},
{32'd4, 32'd5707, 32'd124, -32'd4553},
{-32'd5628, 32'd4974, -32'd8751, -32'd916},
{32'd2348, -32'd11693, 32'd7681, 32'd11470},
{-32'd3136, -32'd2711, 32'd2543, 32'd10408},
{32'd6369, -32'd846, 32'd12364, -32'd2365},
{-32'd6464, -32'd4310, -32'd9346, 32'd8567},
{-32'd13710, -32'd1809, 32'd3748, -32'd7083},
{-32'd5378, -32'd492, 32'd1030, 32'd1062},
{32'd3353, -32'd9100, -32'd1524, -32'd7835},
{-32'd10343, 32'd2192, -32'd3005, 32'd2757},
{-32'd13110, -32'd14135, -32'd1535, 32'd7972},
{-32'd515, -32'd7732, -32'd8161, -32'd3853},
{-32'd1200, -32'd2665, 32'd6782, 32'd5914},
{-32'd1559, 32'd16445, -32'd1192, -32'd1595},
{-32'd9752, -32'd10491, -32'd12017, -32'd848},
{-32'd4583, 32'd934, 32'd8854, 32'd2789},
{-32'd8173, -32'd5357, 32'd2425, -32'd3593},
{32'd1756, -32'd5317, -32'd476, 32'd6275},
{32'd9106, -32'd3775, -32'd4436, 32'd8044},
{-32'd3586, 32'd7244, -32'd934, -32'd1760},
{-32'd5298, -32'd5969, 32'd5129, 32'd3522},
{-32'd6904, -32'd1752, 32'd8235, -32'd5577},
{32'd13135, 32'd6640, 32'd9314, 32'd9329},
{32'd3468, 32'd1204, 32'd7862, 32'd4305},
{-32'd1033, 32'd9710, 32'd9777, 32'd2122},
{32'd3743, 32'd8061, -32'd2468, -32'd8490},
{32'd3018, 32'd9542, -32'd4256, -32'd6932},
{-32'd4393, -32'd2814, -32'd1576, -32'd4362},
{-32'd9454, 32'd7138, -32'd11630, -32'd6677},
{-32'd2344, -32'd3235, -32'd939, -32'd1290},
{32'd2932, 32'd15082, -32'd4247, 32'd3378},
{-32'd3376, 32'd4424, 32'd4775, 32'd769},
{32'd6083, 32'd4692, 32'd5261, 32'd2109},
{-32'd7590, -32'd7933, 32'd2832, 32'd340},
{-32'd45, -32'd1026, -32'd2433, -32'd1953},
{32'd8132, 32'd9167, -32'd7253, 32'd2556},
{32'd16268, 32'd9773, 32'd9186, -32'd1341},
{32'd3318, 32'd15307, 32'd7184, -32'd5165},
{-32'd1984, -32'd3201, 32'd6, -32'd3508},
{-32'd2093, 32'd2348, 32'd7867, -32'd3920},
{-32'd3651, 32'd3619, 32'd5741, 32'd1917},
{-32'd1861, 32'd9313, 32'd5621, -32'd3430},
{32'd6921, 32'd12436, 32'd3607, 32'd3260},
{32'd6118, -32'd3148, 32'd10248, 32'd8122},
{-32'd6960, 32'd2375, 32'd3371, -32'd552},
{-32'd493, 32'd1902, -32'd1841, 32'd1461},
{32'd3262, 32'd4110, -32'd8275, -32'd15243},
{-32'd1463, -32'd16988, -32'd10777, -32'd9769},
{-32'd4154, -32'd10253, 32'd3156, 32'd68},
{-32'd3482, 32'd2689, 32'd2754, -32'd4108},
{-32'd9709, -32'd13708, -32'd4731, -32'd6100},
{32'd5155, 32'd3239, 32'd5164, 32'd4676},
{-32'd11088, -32'd17703, 32'd3343, 32'd5073},
{-32'd10971, 32'd240, 32'd5366, -32'd2632},
{-32'd2372, 32'd14188, -32'd2694, -32'd2530},
{-32'd5301, 32'd164, 32'd2448, 32'd2657},
{32'd2929, 32'd791, 32'd6630, -32'd6322},
{-32'd7342, -32'd761, 32'd3846, 32'd4038},
{-32'd2261, -32'd8951, -32'd3369, -32'd9230},
{32'd10601, -32'd4365, -32'd19473, 32'd66},
{-32'd4488, -32'd420, -32'd13062, 32'd5243},
{32'd99, -32'd4547, 32'd4629, -32'd4897},
{32'd1728, -32'd1640, -32'd12203, 32'd3983},
{32'd145, -32'd7126, 32'd1428, 32'd3310},
{-32'd1357, 32'd6859, 32'd9590, -32'd529},
{32'd6294, -32'd5493, 32'd2574, 32'd1227},
{32'd1587, 32'd4430, -32'd2879, -32'd751},
{-32'd1928, -32'd1070, -32'd4067, -32'd255},
{32'd7890, -32'd5864, -32'd653, 32'd7481},
{-32'd6997, 32'd4000, -32'd7582, 32'd8568},
{-32'd8659, -32'd9947, -32'd12453, -32'd17},
{-32'd13698, -32'd2477, -32'd1052, -32'd2052},
{-32'd7207, 32'd5798, -32'd10042, 32'd1325},
{-32'd5554, -32'd4271, -32'd5490, -32'd1335},
{-32'd7211, 32'd8304, -32'd4188, -32'd5900},
{-32'd11388, 32'd12288, 32'd9977, -32'd7745},
{32'd1615, 32'd4454, 32'd1614, 32'd5637},
{32'd3867, -32'd6826, 32'd9478, -32'd10571},
{-32'd1546, 32'd13914, 32'd1303, 32'd6921},
{-32'd5199, -32'd732, -32'd2858, -32'd7798},
{32'd3826, -32'd15229, -32'd3148, -32'd3492},
{32'd2167, 32'd2983, -32'd8078, -32'd2394},
{32'd3589, -32'd979, 32'd6920, -32'd3928},
{32'd2887, 32'd3145, 32'd171, 32'd9506},
{32'd12049, -32'd6050, 32'd6696, -32'd5640},
{32'd5522, 32'd15320, -32'd529, 32'd9521},
{-32'd4236, 32'd978, 32'd9147, -32'd5066},
{32'd5922, 32'd2339, 32'd1557, -32'd1933},
{32'd5800, 32'd5051, -32'd2603, -32'd825},
{32'd4457, -32'd3542, 32'd1959, 32'd3061},
{32'd3965, 32'd5285, -32'd4162, -32'd5414},
{-32'd4756, 32'd7837, 32'd2596, 32'd3095},
{-32'd1652, 32'd1424, -32'd1336, -32'd12516},
{32'd9564, -32'd4783, -32'd13704, -32'd1819},
{-32'd2858, -32'd4031, -32'd4483, 32'd1656},
{-32'd2629, -32'd1674, 32'd7823, 32'd3132},
{32'd4055, 32'd366, 32'd5602, 32'd3083},
{-32'd961, -32'd4849, 32'd8623, -32'd1264},
{32'd6754, -32'd2110, 32'd8360, -32'd1989},
{-32'd493, -32'd8331, 32'd1157, -32'd11454},
{32'd2324, 32'd9635, 32'd4142, 32'd2406},
{32'd3304, 32'd4980, 32'd136, 32'd1756},
{-32'd5828, -32'd4678, -32'd7263, 32'd1126},
{32'd13533, -32'd679, 32'd3623, 32'd4789},
{32'd3602, 32'd1741, 32'd8578, -32'd369},
{32'd1472, -32'd4477, 32'd8434, -32'd419},
{-32'd452, -32'd4517, -32'd6521, -32'd7724},
{-32'd6066, 32'd4198, -32'd3029, 32'd7615},
{32'd4980, 32'd1646, -32'd8300, 32'd5566},
{-32'd6467, 32'd702, -32'd14468, -32'd12700},
{-32'd9244, 32'd110, -32'd3999, -32'd2148},
{32'd3783, -32'd2643, -32'd567, -32'd7163},
{32'd6803, 32'd1821, 32'd3792, 32'd4288},
{-32'd16764, 32'd2072, 32'd2612, 32'd842},
{-32'd7223, -32'd9507, 32'd2781, 32'd1763},
{-32'd12692, 32'd3221, -32'd1809, 32'd11498},
{-32'd484, -32'd2152, 32'd7124, -32'd541},
{-32'd2400, -32'd4501, 32'd3968, 32'd1621},
{32'd5579, 32'd496, -32'd1872, -32'd7375},
{-32'd682, -32'd30, 32'd704, -32'd3628},
{32'd8091, -32'd9069, 32'd14670, 32'd370},
{32'd912, -32'd9837, -32'd4224, -32'd3903},
{32'd11291, -32'd2398, 32'd258, -32'd6614},
{32'd6347, 32'd13923, 32'd5501, 32'd4270},
{-32'd9976, 32'd2901, -32'd9820, -32'd4661},
{32'd6116, -32'd9080, -32'd5720, 32'd2726},
{32'd117, 32'd1257, -32'd7129, -32'd7055},
{32'd1881, -32'd752, 32'd8927, -32'd89},
{-32'd107, -32'd2352, 32'd8682, 32'd2425},
{32'd6467, -32'd9589, -32'd1294, 32'd5535},
{-32'd10786, 32'd9231, -32'd1545, 32'd9596},
{32'd4246, -32'd4393, -32'd695, 32'd3331},
{32'd18, -32'd4351, 32'd3033, 32'd6144},
{32'd657, 32'd4979, -32'd11608, -32'd18},
{32'd6249, -32'd7514, 32'd76, -32'd406},
{-32'd1075, 32'd6714, -32'd1321, -32'd4641},
{-32'd2208, 32'd8612, -32'd1633, -32'd2662},
{-32'd1126, -32'd431, -32'd7969, -32'd2824},
{32'd2477, -32'd4016, 32'd6285, -32'd5489},
{-32'd3545, 32'd16180, 32'd8425, -32'd2742},
{32'd1319, 32'd6582, 32'd4379, -32'd650},
{32'd5008, -32'd5918, 32'd7498, 32'd7376},
{-32'd2356, -32'd2451, 32'd3626, 32'd526},
{-32'd10029, -32'd903, 32'd12368, 32'd4082},
{-32'd1050, -32'd12701, 32'd10895, -32'd3015},
{-32'd8074, -32'd2502, 32'd2864, 32'd4128},
{32'd594, 32'd1534, -32'd3473, -32'd1842},
{32'd1360, -32'd3152, -32'd4661, 32'd6023},
{32'd3012, -32'd9108, 32'd3311, 32'd3333},
{32'd509, -32'd4423, 32'd5437, 32'd7622},
{32'd1681, 32'd7037, -32'd925, 32'd602},
{32'd594, -32'd1033, 32'd3809, -32'd7306},
{32'd2910, 32'd5705, 32'd1601, 32'd1905},
{-32'd2650, 32'd2400, 32'd3224, 32'd651},
{32'd1527, -32'd1198, 32'd2554, -32'd867},
{32'd4937, 32'd5898, 32'd4218, 32'd6935},
{-32'd5362, 32'd2950, -32'd552, -32'd4319},
{32'd2115, 32'd733, 32'd4098, -32'd6328},
{-32'd7757, 32'd5285, -32'd2504, -32'd406},
{-32'd6799, 32'd12795, 32'd7179, -32'd5346},
{32'd3617, 32'd7109, -32'd1421, -32'd1987},
{32'd2287, 32'd6260, 32'd5519, 32'd5097},
{-32'd7201, -32'd13394, 32'd9353, -32'd12588},
{32'd1291, 32'd4339, 32'd7790, -32'd5581},
{-32'd3910, -32'd8597, -32'd1115, -32'd1066},
{32'd1895, -32'd326, 32'd387, 32'd3709},
{32'd751, 32'd177, -32'd2606, -32'd6288},
{-32'd4478, -32'd11462, 32'd5462, 32'd2043},
{32'd8943, 32'd1618, -32'd7142, 32'd2150},
{32'd2856, -32'd1891, 32'd4279, 32'd7383},
{32'd1856, 32'd2482, 32'd4091, 32'd10843},
{32'd1445, -32'd2034, -32'd1534, 32'd2582},
{-32'd3197, -32'd8769, -32'd8268, -32'd5788},
{-32'd6302, -32'd7486, -32'd8552, -32'd1389},
{-32'd8801, 32'd5879, 32'd3035, 32'd2668},
{32'd4329, 32'd1289, 32'd6738, 32'd567},
{32'd10671, 32'd7510, -32'd2395, 32'd1873},
{-32'd106, 32'd2517, 32'd1410, 32'd1490},
{-32'd8618, 32'd6144, -32'd11161, 32'd982}
},
{{32'd8031, 32'd887, -32'd746, 32'd11502},
{32'd5240, -32'd8520, -32'd797, 32'd4647},
{-32'd7845, 32'd4333, 32'd10069, 32'd6671},
{-32'd542, -32'd529, -32'd3180, 32'd4454},
{32'd6579, 32'd8693, -32'd595, 32'd2362},
{32'd1827, 32'd3613, -32'd8430, 32'd3466},
{-32'd5226, 32'd12734, 32'd4245, 32'd2679},
{32'd104, 32'd1726, -32'd20452, 32'd5893},
{-32'd5144, 32'd1646, -32'd5169, 32'd8516},
{32'd9648, 32'd11653, -32'd1006, -32'd2865},
{32'd7273, -32'd5742, -32'd4760, -32'd442},
{32'd13679, -32'd8840, 32'd6051, -32'd4796},
{-32'd4975, 32'd3749, 32'd5831, -32'd4653},
{32'd7473, -32'd6569, 32'd165, -32'd6021},
{-32'd5174, 32'd3515, -32'd6922, -32'd5447},
{32'd2294, 32'd1480, 32'd4255, -32'd6429},
{32'd6656, -32'd1552, 32'd4956, 32'd6329},
{-32'd7965, 32'd2014, 32'd182, 32'd7046},
{32'd4186, -32'd3676, -32'd12762, -32'd4455},
{32'd7830, 32'd2467, -32'd5176, 32'd6631},
{32'd6683, -32'd2838, -32'd4203, -32'd3058},
{-32'd13369, -32'd4188, -32'd5067, 32'd6993},
{-32'd1710, -32'd2003, -32'd12107, -32'd3697},
{-32'd56, 32'd10191, -32'd4706, -32'd4248},
{32'd12320, 32'd2019, -32'd2997, -32'd3838},
{-32'd6127, -32'd9307, 32'd15031, 32'd4256},
{-32'd4674, -32'd2576, -32'd5960, -32'd2134},
{32'd1747, 32'd6216, 32'd399, 32'd2800},
{32'd6570, 32'd1122, 32'd17778, 32'd4085},
{-32'd13701, 32'd3944, 32'd1872, -32'd11345},
{-32'd4639, 32'd5266, -32'd4168, 32'd4911},
{-32'd3697, -32'd11558, 32'd4559, 32'd2915},
{32'd6903, 32'd7993, -32'd4949, 32'd1264},
{32'd1406, -32'd8040, 32'd6184, -32'd7074},
{32'd1891, 32'd5478, 32'd4737, -32'd2607},
{-32'd7261, -32'd8219, -32'd2457, 32'd8362},
{-32'd6689, 32'd1027, 32'd7129, 32'd9557},
{32'd12769, -32'd10062, 32'd11079, -32'd7948},
{32'd4990, 32'd12500, 32'd3735, -32'd11296},
{-32'd2145, 32'd734, 32'd6466, -32'd6481},
{32'd2261, 32'd10187, 32'd8982, 32'd3587},
{32'd3708, 32'd6510, -32'd885, -32'd3962},
{-32'd8935, -32'd3776, 32'd12146, -32'd6172},
{32'd3004, -32'd5533, -32'd5557, -32'd4560},
{-32'd530, -32'd6390, -32'd9463, -32'd4173},
{32'd4946, -32'd4558, 32'd8121, -32'd10548},
{32'd11903, -32'd4458, -32'd182, 32'd9013},
{32'd8702, -32'd14370, -32'd6832, -32'd978},
{-32'd3779, 32'd7228, -32'd6807, 32'd4936},
{-32'd613, -32'd1547, -32'd1967, -32'd4049},
{32'd333, 32'd3711, 32'd4261, 32'd2483},
{-32'd3584, 32'd1852, -32'd2267, -32'd13509},
{-32'd5857, 32'd905, -32'd1763, 32'd2774},
{-32'd3942, -32'd3513, 32'd3577, 32'd8837},
{32'd9790, 32'd12204, -32'd312, 32'd985},
{32'd8920, 32'd5669, -32'd6509, 32'd16789},
{32'd6950, 32'd13301, 32'd2052, 32'd4138},
{32'd734, 32'd980, -32'd10553, 32'd2652},
{-32'd6432, -32'd5077, -32'd7045, 32'd3977},
{-32'd12724, -32'd5337, -32'd5474, 32'd3963},
{-32'd11268, -32'd3492, 32'd223, 32'd8797},
{-32'd4234, 32'd12639, 32'd15749, -32'd816},
{-32'd17274, 32'd2959, -32'd1541, 32'd216},
{-32'd9643, -32'd7422, 32'd3018, 32'd6914},
{32'd6704, -32'd2237, -32'd7260, -32'd9645},
{32'd10436, -32'd695, -32'd6265, 32'd419},
{32'd6360, -32'd6210, 32'd6473, -32'd6093},
{-32'd12463, 32'd7182, 32'd339, 32'd4278},
{-32'd1577, -32'd103, -32'd8348, -32'd11701},
{-32'd1459, 32'd2194, 32'd677, 32'd7846},
{32'd2440, 32'd3904, -32'd7330, 32'd7236},
{32'd8225, 32'd3042, 32'd4559, 32'd7769},
{32'd281, 32'd3723, 32'd2965, 32'd234},
{32'd15002, 32'd5080, 32'd4565, 32'd2227},
{-32'd1580, -32'd1305, 32'd1099, 32'd5877},
{-32'd9, 32'd1502, 32'd6179, -32'd3047},
{-32'd756, -32'd1244, -32'd4824, -32'd11206},
{-32'd7888, -32'd12427, -32'd10919, -32'd4222},
{-32'd1685, 32'd2097, 32'd10647, 32'd1912},
{-32'd1712, -32'd265, 32'd4295, 32'd246},
{-32'd728, -32'd5177, -32'd15894, -32'd4879},
{32'd207, -32'd984, -32'd4784, -32'd7176},
{32'd10381, 32'd4613, 32'd668, 32'd2642},
{-32'd1252, -32'd192, 32'd11196, 32'd7826},
{-32'd12226, -32'd7488, 32'd2939, -32'd757},
{32'd1206, 32'd11053, 32'd12800, 32'd1858},
{-32'd6225, 32'd8840, 32'd6806, -32'd404},
{-32'd285, -32'd7589, -32'd5208, 32'd885},
{32'd14265, 32'd1782, -32'd3976, -32'd3945},
{32'd2640, -32'd7829, -32'd11920, -32'd5810},
{32'd9710, 32'd4144, -32'd635, -32'd4003},
{-32'd1209, 32'd1179, -32'd2090, 32'd750},
{32'd11387, -32'd3463, -32'd15924, 32'd471},
{-32'd442, 32'd11735, 32'd13590, -32'd2022},
{32'd11082, 32'd6769, 32'd9714, 32'd4724},
{-32'd9925, -32'd10515, -32'd5918, -32'd3029},
{32'd8634, 32'd3550, 32'd3354, -32'd88},
{-32'd7473, 32'd6145, -32'd8702, 32'd3040},
{-32'd8416, 32'd4487, 32'd18667, 32'd4466},
{32'd1516, 32'd4403, -32'd6128, -32'd664},
{-32'd5443, -32'd5182, 32'd5115, -32'd4514},
{32'd817, -32'd1154, 32'd6300, 32'd482},
{32'd10001, 32'd9628, 32'd10635, 32'd89},
{32'd3964, -32'd5857, -32'd9293, -32'd11604},
{-32'd1333, 32'd931, 32'd10272, -32'd5778},
{-32'd1099, -32'd168, 32'd3415, 32'd5629},
{32'd8293, -32'd2406, 32'd11524, -32'd2150},
{32'd8693, -32'd6139, 32'd2490, -32'd10933},
{32'd661, 32'd6961, -32'd3956, -32'd3761},
{-32'd16389, -32'd5007, 32'd10962, 32'd6687},
{32'd8127, 32'd4470, -32'd8806, 32'd2678},
{-32'd2954, 32'd2701, 32'd10582, -32'd7979},
{-32'd2970, -32'd4835, 32'd16604, -32'd554},
{-32'd8140, 32'd2583, 32'd1225, 32'd3808},
{32'd7132, 32'd8763, -32'd1046, -32'd5727},
{-32'd16477, -32'd4200, -32'd659, 32'd1061},
{-32'd1270, -32'd10046, 32'd14467, 32'd6632},
{-32'd3312, -32'd5052, -32'd4133, -32'd5822},
{32'd12594, -32'd7816, -32'd1941, 32'd3271},
{32'd7624, 32'd2623, -32'd1424, 32'd2789},
{-32'd3802, -32'd5726, -32'd6044, -32'd10511},
{-32'd3100, 32'd1544, -32'd3885, 32'd3966},
{32'd3418, -32'd1072, -32'd10371, -32'd3675},
{-32'd1775, 32'd3176, 32'd5735, 32'd5308},
{32'd417, 32'd2082, -32'd3490, 32'd611},
{-32'd3674, 32'd21427, 32'd8590, 32'd5506},
{-32'd4417, -32'd858, -32'd12562, 32'd5437},
{-32'd6275, -32'd4899, -32'd1689, 32'd2051},
{32'd354, -32'd2939, 32'd411, 32'd6732},
{32'd7325, -32'd13642, 32'd2352, 32'd4507},
{32'd2772, 32'd1702, -32'd7844, 32'd6669},
{32'd7709, -32'd1694, -32'd3993, -32'd6291},
{-32'd8241, 32'd5219, -32'd4556, 32'd4797},
{32'd8128, 32'd10756, 32'd10147, 32'd9807},
{-32'd7109, 32'd1625, -32'd18231, 32'd8806},
{32'd13001, 32'd8428, -32'd8863, -32'd1702},
{32'd3292, 32'd3559, -32'd1695, 32'd3173},
{-32'd17416, -32'd786, -32'd5001, 32'd2712},
{32'd8480, -32'd10137, -32'd487, -32'd8552},
{32'd2498, -32'd230, -32'd3827, 32'd4458},
{-32'd127, -32'd464, -32'd7399, -32'd9765},
{32'd4834, 32'd1160, 32'd7974, 32'd6698},
{32'd4276, -32'd23356, -32'd1597, -32'd9876},
{32'd5037, -32'd3335, 32'd4998, 32'd4139},
{-32'd3712, 32'd3155, 32'd4411, 32'd2570},
{32'd929, 32'd5127, -32'd3413, -32'd2920},
{-32'd2050, 32'd3314, 32'd4965, 32'd1321},
{-32'd1636, -32'd324, 32'd7954, 32'd6291},
{32'd2841, 32'd6285, -32'd1692, -32'd633},
{32'd2393, -32'd162, -32'd12021, -32'd2061},
{32'd5009, 32'd2690, 32'd3485, 32'd3414},
{32'd961, -32'd795, 32'd5635, -32'd4432},
{32'd43, 32'd2519, 32'd1798, -32'd3941},
{-32'd5555, 32'd759, 32'd2153, 32'd1154},
{-32'd11385, -32'd3255, 32'd1488, 32'd2110},
{32'd3346, 32'd13351, 32'd3260, 32'd6880},
{32'd958, -32'd15921, -32'd2030, 32'd12038},
{32'd10659, -32'd4307, -32'd502, -32'd3533},
{-32'd2048, 32'd1181, -32'd5933, -32'd8378},
{-32'd10366, -32'd2934, 32'd1568, 32'd6604},
{-32'd3508, -32'd7920, -32'd13618, -32'd1906},
{-32'd2385, 32'd9823, -32'd4501, 32'd4708},
{-32'd8610, 32'd825, 32'd5304, 32'd7731},
{32'd5364, 32'd3436, 32'd11064, 32'd2639},
{32'd8146, -32'd2580, 32'd6978, 32'd3157},
{-32'd2722, -32'd3816, 32'd2532, -32'd16140},
{-32'd6044, 32'd205, 32'd2362, -32'd2340},
{32'd5556, 32'd2153, -32'd2474, 32'd2691},
{-32'd10648, -32'd246, 32'd10387, -32'd2618},
{-32'd13171, -32'd5883, 32'd53, 32'd5327},
{-32'd10274, -32'd9825, -32'd2258, -32'd1651},
{32'd4384, 32'd1636, -32'd20064, 32'd8472},
{32'd729, -32'd3674, 32'd8106, 32'd3775},
{-32'd2499, 32'd3704, 32'd507, -32'd4024},
{32'd8767, -32'd13391, -32'd8897, 32'd10013},
{32'd3970, 32'd6269, -32'd741, -32'd492},
{-32'd2260, -32'd96, 32'd1531, 32'd3049},
{32'd1366, -32'd8248, 32'd8880, 32'd12929},
{32'd20009, 32'd4373, 32'd10269, 32'd3312},
{32'd2537, 32'd2071, -32'd5556, 32'd5821},
{-32'd275, -32'd8263, 32'd619, -32'd8535},
{32'd5304, -32'd3707, -32'd761, -32'd11275},
{-32'd7486, -32'd3793, -32'd846, -32'd646},
{-32'd6764, 32'd2358, -32'd4483, -32'd15410},
{-32'd11398, 32'd6070, -32'd2791, 32'd5619},
{32'd2169, 32'd120, -32'd5147, 32'd4572},
{32'd1782, 32'd2847, -32'd899, 32'd5880},
{32'd1685, -32'd6938, 32'd8033, 32'd2392},
{32'd10277, -32'd3851, -32'd2476, -32'd9624},
{32'd2638, -32'd1635, -32'd4305, -32'd1653},
{-32'd8859, 32'd1954, 32'd5055, 32'd6154},
{32'd1433, -32'd7652, -32'd53, -32'd6050},
{-32'd619, -32'd358, 32'd12626, 32'd1574},
{-32'd676, 32'd4024, -32'd2075, -32'd2905},
{32'd5423, 32'd39, -32'd4870, 32'd650},
{-32'd1384, 32'd7115, -32'd8993, 32'd6312},
{-32'd1082, -32'd9372, 32'd3214, 32'd4466},
{32'd9170, 32'd1786, 32'd401, -32'd6586},
{-32'd2665, 32'd365, -32'd8299, 32'd1387},
{32'd3666, 32'd5302, 32'd5421, 32'd194},
{-32'd4298, -32'd7640, -32'd4867, 32'd2895},
{-32'd7401, 32'd2604, -32'd3594, -32'd1726},
{32'd4763, 32'd7847, 32'd5085, -32'd3659},
{32'd8445, 32'd6939, 32'd3664, 32'd3140},
{32'd16917, -32'd2991, -32'd7350, -32'd13},
{32'd9117, -32'd4758, 32'd12371, 32'd6259},
{-32'd4876, -32'd4802, -32'd20709, 32'd3933},
{32'd12377, -32'd337, 32'd1971, -32'd6479},
{32'd2329, 32'd5942, 32'd609, 32'd5938},
{32'd685, 32'd4697, 32'd3550, 32'd2799},
{-32'd10499, 32'd4351, 32'd12763, -32'd2267},
{32'd3884, -32'd646, 32'd3371, -32'd9507},
{-32'd4214, -32'd3486, -32'd6578, 32'd14581},
{-32'd3178, -32'd17362, 32'd242, -32'd16159},
{-32'd2595, 32'd798, -32'd2978, -32'd304},
{-32'd10124, 32'd2603, -32'd11205, -32'd4931},
{-32'd8422, -32'd5265, 32'd4198, -32'd2742},
{32'd9508, 32'd1306, -32'd2072, -32'd9033},
{-32'd332, 32'd4095, 32'd12021, 32'd1864},
{32'd2474, 32'd3633, 32'd2509, 32'd663},
{32'd2206, 32'd5910, -32'd1237, -32'd2509},
{-32'd17980, -32'd4047, 32'd1976, -32'd892},
{-32'd2021, 32'd8468, 32'd1595, -32'd368},
{32'd1596, -32'd9017, 32'd432, 32'd5678},
{32'd5683, 32'd733, 32'd4286, -32'd1684},
{32'd4322, -32'd12027, 32'd14843, -32'd1414},
{32'd1871, -32'd14568, -32'd17863, -32'd2478},
{-32'd8416, 32'd298, -32'd20908, -32'd3607},
{32'd9689, -32'd9624, -32'd1268, 32'd5169},
{32'd2412, 32'd5888, 32'd6699, 32'd5448},
{-32'd8056, -32'd3256, -32'd4509, -32'd1358},
{32'd1854, -32'd822, 32'd4670, 32'd1873},
{-32'd7159, -32'd5030, 32'd710, -32'd1992},
{-32'd3388, 32'd9217, -32'd12001, -32'd1301},
{32'd2893, -32'd2404, -32'd6482, 32'd1432},
{-32'd9740, -32'd2221, -32'd773, 32'd10882},
{32'd9750, -32'd2394, -32'd1956, -32'd11983},
{-32'd4107, 32'd4099, 32'd10165, -32'd2715},
{-32'd1360, 32'd1613, -32'd3419, 32'd2726},
{-32'd873, -32'd244, -32'd11292, -32'd3544},
{32'd1038, 32'd12536, 32'd6668, 32'd5356},
{-32'd470, -32'd3263, -32'd3328, -32'd864},
{-32'd3982, -32'd279, -32'd5383, 32'd4131},
{-32'd5281, 32'd2649, 32'd2958, -32'd10849},
{32'd7594, 32'd8786, 32'd1085, -32'd1007},
{32'd2405, -32'd2936, -32'd12063, -32'd247},
{-32'd1074, 32'd10737, 32'd6123, -32'd1687},
{32'd2533, 32'd1006, -32'd9410, 32'd11220},
{32'd11022, -32'd8230, -32'd9010, 32'd4372},
{32'd4072, 32'd2766, 32'd15745, -32'd704},
{-32'd7258, -32'd1510, -32'd15022, -32'd13215},
{-32'd5573, 32'd1856, -32'd9482, -32'd4666},
{32'd4671, 32'd5607, -32'd7968, 32'd3206},
{-32'd2213, -32'd6841, -32'd7274, -32'd8367},
{-32'd2394, -32'd5985, -32'd625, -32'd12701},
{-32'd2652, -32'd1726, 32'd15610, 32'd5985},
{32'd2830, 32'd4636, 32'd898, -32'd3714},
{32'd1963, 32'd4940, -32'd5433, -32'd2765},
{32'd2840, -32'd6632, -32'd15025, -32'd4119},
{32'd2304, 32'd1585, 32'd10391, -32'd3662},
{-32'd163, -32'd4, 32'd882, 32'd1929},
{32'd9855, 32'd931, 32'd13362, 32'd5639},
{-32'd10451, -32'd1434, 32'd5741, -32'd7638},
{32'd1186, -32'd568, 32'd250, -32'd1338},
{32'd2420, -32'd10109, -32'd3643, -32'd1816},
{32'd2184, -32'd4722, 32'd7733, 32'd667},
{32'd1554, 32'd6115, 32'd3577, 32'd168},
{-32'd15562, -32'd3901, 32'd11450, 32'd8266},
{32'd6420, -32'd5200, -32'd5609, 32'd4131},
{-32'd14113, 32'd3096, 32'd2990, 32'd3145},
{32'd5146, -32'd16201, -32'd710, -32'd5436},
{32'd3429, -32'd2534, -32'd8415, 32'd7520},
{32'd3175, -32'd2108, 32'd8345, 32'd6363},
{-32'd11774, -32'd7120, -32'd7057, 32'd3961},
{32'd7620, 32'd2092, -32'd6309, 32'd1590},
{32'd6595, -32'd14457, 32'd5999, 32'd7305},
{32'd5384, 32'd11104, -32'd740, -32'd2444},
{-32'd4012, 32'd3965, 32'd2274, -32'd5181},
{-32'd3523, -32'd2835, -32'd981, 32'd3176},
{32'd6570, 32'd6685, 32'd6517, -32'd1189},
{32'd12298, -32'd2410, -32'd10248, 32'd5602},
{32'd1233, -32'd7864, 32'd6949, 32'd2619},
{32'd6972, -32'd7858, 32'd12864, 32'd10752},
{-32'd909, -32'd2306, -32'd5542, 32'd276},
{-32'd4105, -32'd6061, 32'd3855, -32'd5455},
{-32'd3617, 32'd8083, -32'd1646, -32'd3085},
{-32'd217, 32'd5217, -32'd10258, 32'd4900},
{-32'd18350, 32'd4025, -32'd1785, -32'd5767},
{32'd1130, -32'd208, 32'd2133, 32'd8124},
{-32'd341, 32'd9694, 32'd1539, 32'd4948},
{32'd319, 32'd2383, 32'd927, 32'd5777},
{-32'd246, 32'd6116, 32'd1356, -32'd4680},
{32'd1503, -32'd3277, 32'd4180, 32'd5705},
{32'd785, 32'd989, 32'd4308, -32'd11625},
{32'd2497, -32'd3395, 32'd1609, 32'd474},
{32'd2128, 32'd1222, -32'd7523, -32'd3053},
{-32'd2753, 32'd2839, 32'd9344, -32'd4420},
{-32'd6536, 32'd4806, -32'd6546, 32'd171},
{32'd11374, 32'd3375, -32'd1724, -32'd6195},
{32'd1121, -32'd10372, -32'd13555, 32'd1338}
},
{{-32'd14738, 32'd14684, -32'd895, -32'd1103},
{-32'd11135, -32'd7569, -32'd16089, -32'd4294},
{32'd363, -32'd8376, 32'd4102, 32'd1687},
{32'd12831, 32'd3970, 32'd2893, 32'd3896},
{32'd7747, -32'd2645, -32'd4688, 32'd17614},
{32'd9464, -32'd4389, 32'd2095, -32'd5791},
{-32'd10424, 32'd1789, 32'd12995, 32'd210},
{-32'd3119, 32'd3395, -32'd6958, -32'd1979},
{32'd6675, -32'd2610, 32'd753, 32'd2174},
{32'd2804, 32'd11764, 32'd7147, 32'd11479},
{-32'd3114, -32'd7853, -32'd10382, 32'd5227},
{-32'd9280, 32'd2459, -32'd4768, -32'd280},
{-32'd4562, 32'd5885, -32'd8525, 32'd10454},
{32'd5620, -32'd5624, -32'd3888, -32'd4807},
{-32'd1319, 32'd3268, 32'd366, -32'd5824},
{-32'd7962, 32'd881, 32'd6714, -32'd8536},
{-32'd1695, 32'd16920, 32'd10317, -32'd3554},
{32'd497, -32'd4500, -32'd5435, -32'd13867},
{32'd429, 32'd7985, 32'd8793, 32'd14784},
{32'd2171, 32'd3235, 32'd678, 32'd1662},
{-32'd2736, 32'd5659, 32'd3977, 32'd5666},
{-32'd5070, -32'd15540, 32'd1168, -32'd11041},
{32'd832, -32'd58, 32'd3611, -32'd7277},
{32'd2072, -32'd11095, 32'd874, -32'd1416},
{32'd19021, 32'd9331, -32'd1189, 32'd8774},
{32'd11218, 32'd2007, 32'd9058, -32'd1435},
{-32'd6418, -32'd2258, 32'd3387, -32'd2314},
{-32'd6727, 32'd9798, -32'd6170, 32'd1737},
{-32'd8758, 32'd344, 32'd2846, -32'd3688},
{32'd1847, -32'd6408, -32'd5841, 32'd3848},
{-32'd76, 32'd2321, -32'd9636, -32'd2055},
{32'd1763, -32'd12594, -32'd3078, 32'd991},
{32'd8041, 32'd4832, 32'd5016, -32'd2025},
{32'd9500, -32'd8548, -32'd9617, -32'd3627},
{32'd8337, 32'd4737, 32'd7528, 32'd10627},
{-32'd1408, -32'd8782, -32'd4384, 32'd1251},
{-32'd5570, 32'd3862, 32'd261, -32'd7110},
{32'd4587, 32'd4324, -32'd6557, 32'd8075},
{-32'd15681, -32'd5865, 32'd1514, -32'd8094},
{32'd5360, -32'd6159, 32'd2091, -32'd4869},
{-32'd2289, -32'd14682, 32'd3507, -32'd3453},
{-32'd4651, 32'd2897, -32'd11250, 32'd3549},
{-32'd10559, -32'd2556, -32'd3508, 32'd8518},
{-32'd423, 32'd998, 32'd4346, 32'd569},
{32'd8120, -32'd8750, -32'd6905, -32'd5354},
{32'd4719, -32'd213, -32'd3486, 32'd15455},
{32'd1628, -32'd4494, -32'd9029, 32'd14198},
{32'd7816, -32'd830, -32'd5192, 32'd3694},
{32'd1941, -32'd66, 32'd4584, 32'd6015},
{-32'd9291, -32'd4309, -32'd12120, 32'd96},
{-32'd6281, -32'd4369, -32'd2515, 32'd2450},
{32'd6014, 32'd448, -32'd4899, 32'd837},
{-32'd10937, -32'd5382, -32'd417, 32'd5323},
{32'd251, 32'd1009, -32'd4403, 32'd891},
{32'd8353, -32'd3274, 32'd21379, -32'd15817},
{-32'd1988, -32'd448, -32'd12553, -32'd3203},
{-32'd121, 32'd2182, -32'd4042, 32'd7288},
{32'd7986, 32'd257, -32'd9657, 32'd5363},
{-32'd2791, -32'd7468, 32'd4396, 32'd11767},
{-32'd5333, -32'd2018, 32'd1305, -32'd4602},
{32'd228, 32'd3413, 32'd5627, 32'd2872},
{-32'd6355, -32'd17121, -32'd4717, 32'd3579},
{-32'd6837, -32'd8673, -32'd250, 32'd1982},
{-32'd7470, 32'd6232, -32'd2272, -32'd1378},
{32'd8029, 32'd6236, -32'd14155, 32'd9175},
{-32'd10591, 32'd3125, 32'd756, 32'd7032},
{-32'd9725, 32'd8722, 32'd1930, -32'd4216},
{-32'd10794, 32'd30, 32'd3939, -32'd1944},
{-32'd8080, -32'd8921, -32'd12589, -32'd11661},
{-32'd1080, -32'd7544, 32'd9433, -32'd2063},
{-32'd559, 32'd20, -32'd5345, -32'd9549},
{-32'd8420, -32'd5960, -32'd7745, -32'd13602},
{32'd1967, 32'd673, -32'd1581, -32'd13783},
{-32'd11922, -32'd2953, -32'd2612, -32'd9497},
{32'd11145, -32'd3953, 32'd9293, 32'd459},
{32'd6463, -32'd5748, -32'd5193, -32'd6210},
{32'd9527, -32'd8220, -32'd10078, 32'd3432},
{-32'd4342, 32'd6570, 32'd2914, -32'd845},
{32'd775, 32'd11558, 32'd823, -32'd1046},
{-32'd228, -32'd7441, 32'd2142, -32'd3921},
{32'd7994, 32'd7831, 32'd4028, 32'd6668},
{-32'd4585, 32'd11756, -32'd983, 32'd5630},
{-32'd7104, -32'd1364, -32'd2745, 32'd2957},
{-32'd12688, 32'd2463, -32'd450, -32'd6300},
{32'd4407, -32'd13841, -32'd3329, -32'd4283},
{-32'd2486, -32'd1720, 32'd3840, 32'd2066},
{32'd1132, -32'd59, -32'd6802, 32'd5527},
{-32'd9555, -32'd728, -32'd3851, -32'd6170},
{32'd6325, -32'd3092, -32'd14112, 32'd11236},
{-32'd4606, 32'd3153, -32'd879, -32'd7841},
{32'd3040, 32'd7756, -32'd1829, 32'd15265},
{-32'd8284, -32'd3431, -32'd6618, -32'd8357},
{-32'd1543, 32'd2112, -32'd4186, 32'd9325},
{-32'd1361, 32'd2397, 32'd7557, 32'd8444},
{-32'd5115, -32'd2, 32'd4001, 32'd8853},
{32'd1285, -32'd13566, -32'd7876, 32'd752},
{32'd361, 32'd2420, 32'd5616, 32'd14312},
{32'd5030, 32'd2169, 32'd1577, 32'd1429},
{-32'd3193, -32'd11038, 32'd2493, -32'd8379},
{32'd10635, 32'd7042, 32'd2324, 32'd12481},
{-32'd3766, -32'd8389, 32'd12106, 32'd4248},
{-32'd909, -32'd8920, -32'd1779, -32'd5352},
{32'd6995, 32'd628, 32'd13492, 32'd949},
{32'd7040, -32'd906, 32'd1953, 32'd8522},
{32'd2982, 32'd4088, 32'd2076, 32'd4151},
{-32'd5621, -32'd15816, 32'd8550, -32'd4220},
{32'd13090, 32'd1909, -32'd3930, 32'd3104},
{-32'd5662, 32'd1763, -32'd3449, -32'd15103},
{32'd4214, 32'd3367, 32'd12293, 32'd2082},
{-32'd5658, -32'd1823, 32'd2697, 32'd9498},
{-32'd6412, -32'd8154, -32'd5152, -32'd8149},
{32'd829, -32'd1484, -32'd968, 32'd4094},
{-32'd2885, 32'd1121, -32'd10283, 32'd7755},
{-32'd2272, -32'd5174, 32'd545, 32'd11479},
{32'd259, 32'd279, 32'd2777, 32'd7352},
{-32'd15884, 32'd10896, 32'd1444, -32'd11270},
{-32'd6382, -32'd2100, 32'd12596, 32'd361},
{32'd7683, 32'd2997, 32'd10515, -32'd1040},
{32'd8266, -32'd2826, -32'd1214, 32'd6472},
{-32'd10758, 32'd3439, 32'd6420, 32'd5715},
{-32'd1482, 32'd4103, -32'd2008, -32'd5627},
{32'd2566, -32'd10851, -32'd4075, 32'd10379},
{-32'd10611, -32'd8472, 32'd2899, -32'd7057},
{32'd4302, -32'd1509, 32'd6760, 32'd7110},
{32'd471, -32'd7969, 32'd1787, 32'd14076},
{32'd8306, -32'd501, 32'd3528, 32'd1967},
{32'd10302, -32'd2151, 32'd2298, 32'd6926},
{32'd5442, 32'd206, -32'd4303, -32'd6153},
{-32'd3700, -32'd1743, 32'd5761, 32'd8093},
{-32'd1758, 32'd5108, -32'd3835, -32'd7013},
{-32'd18162, 32'd2331, 32'd9000, -32'd1027},
{32'd4782, -32'd9279, -32'd1191, 32'd4220},
{-32'd1860, -32'd11118, 32'd10945, -32'd1872},
{32'd617, -32'd6482, -32'd405, -32'd7090},
{32'd2944, 32'd13026, -32'd12299, 32'd8649},
{-32'd6709, -32'd4656, -32'd11876, -32'd2561},
{32'd8495, -32'd2320, -32'd3140, -32'd2960},
{-32'd7286, -32'd1801, -32'd8791, 32'd14033},
{32'd12907, 32'd13026, 32'd8020, 32'd8030},
{-32'd6760, -32'd10583, 32'd11744, -32'd8888},
{-32'd7259, -32'd4452, 32'd7023, -32'd941},
{32'd1607, -32'd9628, -32'd2323, -32'd13807},
{-32'd8966, 32'd11402, -32'd1783, -32'd13128},
{-32'd6420, -32'd7862, 32'd11239, 32'd6370},
{-32'd3479, -32'd1373, 32'd3814, -32'd1683},
{-32'd1351, 32'd11023, 32'd10438, -32'd1975},
{-32'd8484, 32'd2522, -32'd499, 32'd6019},
{32'd7938, -32'd406, 32'd8355, -32'd160},
{32'd2351, 32'd3514, 32'd3657, 32'd1812},
{-32'd905, -32'd4698, 32'd1953, 32'd5362},
{-32'd66, -32'd1498, -32'd10194, -32'd8744},
{-32'd5051, 32'd6374, -32'd1814, -32'd2625},
{-32'd5898, 32'd1002, 32'd2714, 32'd5636},
{32'd1238, 32'd3110, 32'd2938, 32'd9956},
{32'd869, -32'd7912, -32'd12385, -32'd1048},
{32'd16603, 32'd9179, -32'd2240, -32'd3589},
{-32'd4217, 32'd1991, 32'd10425, 32'd6693},
{32'd7132, -32'd6149, 32'd39, -32'd2692},
{32'd8016, 32'd3390, -32'd1770, -32'd2666},
{-32'd4394, 32'd6157, 32'd1099, 32'd10402},
{32'd3567, -32'd2474, -32'd10866, -32'd5722},
{32'd7459, 32'd466, -32'd2300, -32'd5043},
{-32'd12239, 32'd653, -32'd9936, 32'd6693},
{32'd1099, 32'd7422, -32'd5929, -32'd5014},
{32'd11990, 32'd817, 32'd3112, -32'd4240},
{32'd2595, -32'd1187, -32'd6129, -32'd54},
{32'd602, 32'd10702, 32'd8144, -32'd14388},
{32'd977, -32'd11991, -32'd13720, -32'd14446},
{-32'd10398, 32'd322, -32'd4140, -32'd1768},
{-32'd4744, -32'd1732, -32'd1051, -32'd16647},
{-32'd9616, -32'd12121, -32'd5500, -32'd5246},
{32'd11343, 32'd2676, 32'd22678, 32'd6165},
{32'd7895, 32'd8647, 32'd5868, 32'd10235},
{-32'd1198, 32'd339, -32'd3863, 32'd1283},
{-32'd521, 32'd5837, -32'd5539, 32'd8835},
{-32'd4551, -32'd443, -32'd16341, 32'd747},
{-32'd4771, 32'd9323, 32'd12499, 32'd5360},
{-32'd5607, 32'd7202, -32'd4818, -32'd3901},
{-32'd708, 32'd5661, -32'd3075, 32'd10092},
{-32'd5165, -32'd11962, 32'd4771, -32'd3956},
{-32'd12336, 32'd7327, 32'd3219, -32'd17045},
{32'd1370, -32'd1671, -32'd2498, -32'd2205},
{-32'd3400, -32'd360, -32'd12280, -32'd1299},
{-32'd7256, -32'd7926, -32'd19370, -32'd5666},
{32'd814, -32'd6686, 32'd4277, -32'd6914},
{32'd2914, 32'd7329, -32'd76, 32'd15744},
{-32'd5678, 32'd3731, -32'd2111, -32'd1578},
{32'd5816, -32'd1317, -32'd16272, -32'd9333},
{32'd4908, 32'd11154, -32'd178, -32'd2178},
{32'd6008, -32'd4929, 32'd1703, -32'd1105},
{32'd19001, -32'd1777, -32'd5822, 32'd6406},
{32'd7204, -32'd2393, -32'd2192, -32'd147},
{32'd5034, -32'd1183, -32'd1360, -32'd2751},
{32'd2956, 32'd84, 32'd8845, -32'd1211},
{-32'd8131, 32'd7058, -32'd10566, -32'd13487},
{32'd13787, -32'd1940, 32'd13339, -32'd1800},
{-32'd1533, 32'd388, 32'd8433, 32'd9165},
{-32'd6366, 32'd2310, -32'd4777, -32'd7379},
{-32'd7589, -32'd2299, 32'd259, -32'd6661},
{-32'd4478, 32'd4999, 32'd1253, 32'd2490},
{-32'd1199, -32'd10666, -32'd8456, -32'd6845},
{32'd5696, -32'd5597, 32'd5690, -32'd9777},
{-32'd6549, -32'd4845, -32'd4072, 32'd8300},
{32'd17897, 32'd15252, -32'd6071, 32'd2669},
{32'd6668, -32'd12649, -32'd15456, 32'd3331},
{-32'd3178, -32'd4469, -32'd2658, -32'd7845},
{32'd6180, 32'd8599, 32'd5204, -32'd7380},
{-32'd13008, 32'd979, -32'd10796, -32'd10831},
{-32'd6544, -32'd1058, 32'd6890, -32'd6311},
{-32'd2544, -32'd5435, 32'd5574, 32'd3313},
{32'd1593, -32'd8666, -32'd6453, -32'd8512},
{-32'd5819, 32'd5663, -32'd9719, 32'd2487},
{32'd6805, -32'd12920, -32'd5741, -32'd5251},
{32'd2026, -32'd7165, -32'd4843, -32'd3495},
{32'd4599, -32'd3194, 32'd11039, 32'd5885},
{32'd11383, -32'd664, 32'd9811, -32'd8677},
{32'd2835, 32'd5648, 32'd6497, 32'd1986},
{-32'd4599, 32'd3090, -32'd437, -32'd17863},
{-32'd9400, 32'd4499, 32'd13157, 32'd1778},
{-32'd2293, -32'd8743, -32'd12353, 32'd1958},
{32'd712, 32'd685, -32'd7505, 32'd13670},
{-32'd2760, 32'd4787, 32'd2818, 32'd8193},
{32'd5360, 32'd9686, 32'd7516, 32'd4916},
{32'd7647, -32'd4522, -32'd9944, 32'd877},
{-32'd1824, 32'd2704, 32'd995, 32'd8847},
{32'd1018, -32'd10827, 32'd3835, -32'd3979},
{32'd7504, 32'd5730, -32'd4471, -32'd3271},
{32'd3534, -32'd6677, -32'd6615, -32'd9658},
{-32'd8316, -32'd6768, 32'd7547, 32'd6260},
{-32'd3878, 32'd526, 32'd19428, 32'd2263},
{-32'd9893, 32'd2333, -32'd4317, 32'd2180},
{-32'd8879, -32'd2549, 32'd11110, 32'd1145},
{-32'd7194, 32'd7116, 32'd4663, 32'd1767},
{32'd13914, -32'd3314, -32'd4693, -32'd1333},
{32'd14440, 32'd2274, -32'd5420, 32'd1030},
{32'd6537, -32'd2640, -32'd19147, -32'd8130},
{32'd414, -32'd8579, -32'd14701, -32'd4355},
{-32'd6789, 32'd7003, 32'd6451, 32'd5772},
{32'd12804, -32'd993, 32'd1437, 32'd4996},
{32'd131, -32'd15168, -32'd13446, -32'd5736},
{-32'd14124, -32'd8678, -32'd4500, 32'd4576},
{-32'd81, -32'd3704, -32'd14826, 32'd345},
{-32'd151, -32'd10758, 32'd5647, -32'd13258},
{32'd9253, -32'd10540, 32'd6340, -32'd5659},
{32'd10452, 32'd12804, -32'd430, 32'd2422},
{32'd6866, 32'd11638, -32'd1135, -32'd3864},
{-32'd5652, 32'd729, 32'd7109, -32'd5564},
{32'd8562, -32'd5897, 32'd1194, 32'd5824},
{32'd7061, 32'd725, 32'd3708, -32'd3959},
{-32'd388, 32'd4144, 32'd8708, -32'd4009},
{-32'd3906, 32'd6893, -32'd7537, 32'd3900},
{32'd11202, -32'd968, 32'd9302, 32'd5604},
{32'd17183, 32'd9843, 32'd894, -32'd353},
{-32'd4968, 32'd14122, 32'd6511, 32'd6346},
{-32'd5582, 32'd1792, 32'd8357, -32'd3333},
{-32'd5122, 32'd225, 32'd6495, 32'd15659},
{-32'd4455, 32'd13150, 32'd469, 32'd3865},
{32'd11836, 32'd5766, 32'd10214, 32'd7302},
{-32'd7685, -32'd16, -32'd1648, -32'd5754},
{-32'd2246, 32'd4969, 32'd6363, -32'd6913},
{32'd6958, 32'd14366, 32'd2720, -32'd526},
{32'd8313, 32'd7007, -32'd11395, 32'd6897},
{32'd9505, -32'd20369, -32'd6810, 32'd7330},
{32'd4050, -32'd7831, -32'd14651, -32'd7466},
{32'd7578, 32'd9095, -32'd6567, 32'd6276},
{-32'd5981, -32'd5705, 32'd1114, 32'd6096},
{32'd2938, 32'd8080, 32'd7729, 32'd3758},
{-32'd8391, -32'd14096, -32'd9116, -32'd5505},
{32'd3038, -32'd13235, -32'd298, 32'd8881},
{-32'd217, 32'd512, -32'd6229, 32'd3629},
{-32'd6211, 32'd3443, 32'd7114, 32'd1164},
{32'd2898, -32'd915, 32'd3295, -32'd1575},
{32'd4583, -32'd4974, -32'd6601, -32'd512},
{32'd11171, 32'd1194, -32'd2187, -32'd12706},
{32'd8366, -32'd5494, -32'd845, 32'd2031},
{32'd4565, -32'd4804, -32'd10294, 32'd3746},
{32'd6527, 32'd8339, 32'd5988, 32'd10935},
{-32'd7433, -32'd890, 32'd4422, -32'd1740},
{32'd2700, -32'd8464, -32'd2771, -32'd14496},
{-32'd4424, -32'd9988, 32'd2629, -32'd3834},
{32'd14909, 32'd487, -32'd1580, 32'd1028},
{32'd8072, 32'd3312, -32'd6548, 32'd5475},
{-32'd11020, -32'd4333, -32'd1571, -32'd1818},
{-32'd14869, -32'd5555, -32'd1088, -32'd2751},
{32'd5837, -32'd580, -32'd7489, -32'd9229},
{-32'd9803, -32'd901, -32'd2021, -32'd3627},
{-32'd9885, 32'd10028, 32'd5200, -32'd2063},
{-32'd783, -32'd6092, -32'd554, 32'd192},
{-32'd6101, -32'd2548, -32'd11301, 32'd3707},
{32'd4787, -32'd9460, -32'd8112, -32'd166},
{32'd6975, -32'd1216, 32'd3446, 32'd7707},
{-32'd998, 32'd13718, 32'd48, 32'd4287},
{32'd1747, 32'd6843, 32'd3272, 32'd4177},
{-32'd8313, -32'd10091, -32'd8132, -32'd2330},
{-32'd22712, -32'd2126, -32'd3701, -32'd7395},
{-32'd2158, -32'd10054, -32'd8545, -32'd11830},
{32'd9732, -32'd2769, -32'd4121, -32'd4440},
{32'd1626, -32'd4027, 32'd2115, -32'd3654},
{32'd8982, 32'd1546, 32'd8363, -32'd11616},
{-32'd2640, -32'd2686, 32'd46, 32'd5703}
},
{{32'd2317, 32'd9896, 32'd992, 32'd11227},
{-32'd15237, -32'd6530, -32'd4742, -32'd759},
{32'd6215, 32'd6243, 32'd7347, 32'd8375},
{32'd19399, 32'd3584, 32'd3901, 32'd3554},
{-32'd1206, 32'd5353, 32'd1663, 32'd5819},
{-32'd8324, 32'd8481, -32'd3908, 32'd371},
{32'd1264, 32'd2698, -32'd8757, -32'd9590},
{-32'd10984, 32'd2858, 32'd2554, 32'd583},
{-32'd5432, -32'd1649, -32'd9560, -32'd2971},
{32'd5335, 32'd11185, 32'd2780, 32'd1395},
{-32'd5910, 32'd1894, -32'd4864, 32'd1787},
{-32'd1044, 32'd1598, -32'd2299, -32'd11088},
{-32'd10547, 32'd10652, 32'd2849, -32'd3962},
{-32'd3779, -32'd8431, 32'd118, 32'd6380},
{-32'd6933, -32'd8223, -32'd5725, -32'd6258},
{32'd5553, -32'd1557, -32'd1233, 32'd109},
{-32'd2093, -32'd6325, 32'd3329, 32'd10697},
{32'd3184, 32'd249, 32'd3266, -32'd8441},
{-32'd6292, 32'd3852, -32'd7637, -32'd3436},
{32'd1012, -32'd5262, 32'd810, 32'd2848},
{32'd348, -32'd3741, -32'd131, 32'd636},
{-32'd2791, 32'd341, -32'd2540, 32'd265},
{32'd4893, -32'd4450, -32'd8521, 32'd9628},
{32'd70, 32'd4468, 32'd1072, 32'd6204},
{32'd1227, 32'd5043, 32'd3550, -32'd2597},
{32'd10243, 32'd4659, -32'd8908, 32'd3059},
{32'd1165, 32'd920, -32'd3304, -32'd189},
{-32'd2268, 32'd7684, 32'd2906, -32'd5896},
{-32'd1368, -32'd1046, 32'd2836, 32'd9621},
{-32'd1531, 32'd1063, -32'd4672, -32'd339},
{-32'd5081, 32'd8204, -32'd4144, -32'd4419},
{-32'd1306, -32'd5163, -32'd6480, 32'd6610},
{32'd2072, 32'd2404, -32'd3785, -32'd3279},
{-32'd7228, -32'd2223, 32'd8928, -32'd3029},
{32'd4260, 32'd10466, 32'd3102, -32'd148},
{32'd377, -32'd168, -32'd11900, 32'd3337},
{32'd8622, -32'd6436, 32'd8693, -32'd3189},
{-32'd7340, -32'd4569, -32'd2772, 32'd1193},
{-32'd4512, -32'd1744, -32'd3099, 32'd961},
{32'd4456, -32'd2814, 32'd469, -32'd9788},
{-32'd3517, -32'd8196, -32'd139, -32'd3452},
{32'd6928, 32'd10419, -32'd4579, 32'd533},
{32'd3564, 32'd6768, -32'd2857, -32'd1464},
{-32'd8941, -32'd5946, 32'd1241, -32'd3784},
{-32'd8513, 32'd3785, 32'd6526, 32'd309},
{-32'd9627, -32'd11614, 32'd7437, -32'd3248},
{-32'd7014, 32'd2840, 32'd7505, -32'd1885},
{32'd6846, -32'd4059, 32'd8695, 32'd6338},
{-32'd853, 32'd4201, -32'd3516, 32'd10010},
{-32'd6198, 32'd6264, 32'd3872, -32'd4593},
{32'd2550, -32'd4484, 32'd7648, -32'd2145},
{32'd8418, -32'd5169, 32'd3038, -32'd7135},
{32'd379, 32'd1745, -32'd5692, 32'd4067},
{-32'd17305, -32'd6528, -32'd12372, 32'd14511},
{-32'd4599, -32'd7158, -32'd4245, 32'd1173},
{32'd2678, 32'd668, 32'd5838, 32'd1403},
{-32'd2046, 32'd2453, 32'd9955, 32'd8598},
{32'd898, -32'd5612, -32'd11413, -32'd2264},
{-32'd3824, 32'd2315, 32'd2746, -32'd10663},
{-32'd572, 32'd3205, 32'd7671, -32'd5319},
{-32'd1854, -32'd1380, 32'd8465, 32'd14358},
{32'd5644, -32'd4035, -32'd145, 32'd5310},
{-32'd4075, -32'd1091, -32'd5869, 32'd4652},
{32'd4791, 32'd5495, -32'd3302, -32'd8308},
{-32'd6301, -32'd1790, 32'd12006, -32'd1909},
{-32'd100, 32'd11051, 32'd5330, 32'd7002},
{-32'd11023, 32'd1961, 32'd10073, -32'd15578},
{-32'd3825, -32'd480, -32'd6425, 32'd12232},
{-32'd4755, -32'd134, -32'd1857, 32'd4538},
{-32'd2406, -32'd1126, 32'd1324, 32'd443},
{-32'd2300, -32'd3322, 32'd1614, -32'd5363},
{32'd6162, 32'd5280, 32'd6278, 32'd3317},
{32'd6184, -32'd2791, -32'd5766, -32'd8023},
{-32'd6948, -32'd2456, 32'd2211, -32'd13352},
{32'd416, 32'd2743, -32'd273, 32'd3397},
{-32'd7618, 32'd10297, 32'd9905, -32'd5337},
{-32'd9217, -32'd4175, 32'd4411, -32'd9472},
{-32'd3840, -32'd4082, -32'd6948, -32'd106},
{32'd5889, 32'd3922, 32'd7575, -32'd3692},
{32'd2371, 32'd5229, 32'd5963, 32'd3437},
{32'd13653, -32'd420, -32'd3016, -32'd1789},
{32'd4986, -32'd2830, 32'd1280, -32'd730},
{32'd1696, 32'd2770, -32'd1842, -32'd3978},
{-32'd3677, -32'd1785, -32'd1278, 32'd1481},
{32'd9392, -32'd637, -32'd89, -32'd1750},
{32'd7975, -32'd60, -32'd14789, -32'd538},
{-32'd3584, 32'd8185, 32'd6700, 32'd5603},
{-32'd5575, 32'd293, -32'd453, 32'd4276},
{-32'd7360, 32'd3987, 32'd12824, 32'd5328},
{-32'd4288, -32'd1608, 32'd671, 32'd3608},
{-32'd1651, 32'd3745, 32'd5194, 32'd2754},
{32'd2207, -32'd5699, -32'd4822, 32'd177},
{32'd5434, 32'd4681, 32'd2435, 32'd13391},
{32'd1847, -32'd1229, 32'd7866, 32'd7631},
{32'd2044, 32'd3580, -32'd1168, -32'd6783},
{-32'd13696, 32'd7380, -32'd2964, 32'd9220},
{32'd4491, 32'd7826, 32'd13442, 32'd2191},
{-32'd3985, 32'd3551, -32'd1451, -32'd2015},
{32'd8495, -32'd7, -32'd6353, 32'd5843},
{32'd9507, 32'd5724, 32'd3190, -32'd62},
{-32'd6754, 32'd1250, 32'd1534, -32'd4968},
{-32'd2558, 32'd1514, -32'd2998, -32'd2385},
{32'd1743, 32'd1712, 32'd93, -32'd2785},
{-32'd4306, -32'd4210, 32'd5065, 32'd4216},
{32'd6761, 32'd5990, 32'd3059, -32'd4408},
{-32'd4773, 32'd695, -32'd12701, -32'd2762},
{-32'd13014, 32'd5033, -32'd8103, 32'd1689},
{32'd13574, -32'd855, 32'd9442, 32'd10560},
{32'd3798, 32'd3249, 32'd7897, 32'd5960},
{-32'd3552, -32'd15, 32'd603, -32'd3091},
{32'd2701, -32'd12811, 32'd8557, 32'd5100},
{-32'd1356, 32'd1881, 32'd1569, -32'd3584},
{-32'd45, -32'd1365, 32'd7423, 32'd17424},
{-32'd863, 32'd7309, 32'd9383, 32'd7},
{-32'd4229, 32'd7582, -32'd8129, 32'd4450},
{32'd2982, -32'd6283, -32'd3714, -32'd2402},
{32'd9306, 32'd6227, 32'd4436, 32'd3178},
{-32'd4052, 32'd2496, -32'd6924, 32'd3162},
{-32'd1264, -32'd3640, -32'd10629, -32'd4320},
{32'd13848, 32'd8434, -32'd12828, -32'd27},
{32'd7443, 32'd4128, -32'd2020, 32'd10194},
{-32'd1076, -32'd2769, -32'd417, -32'd4531},
{-32'd14564, -32'd5884, 32'd2413, 32'd610},
{-32'd3348, 32'd722, -32'd2299, -32'd2174},
{32'd12030, 32'd3148, 32'd1767, -32'd9008},
{-32'd2678, -32'd7478, 32'd1871, -32'd9650},
{-32'd1654, 32'd845, -32'd8652, -32'd11660},
{-32'd6451, 32'd1432, -32'd6043, 32'd3692},
{-32'd9362, 32'd10064, -32'd6457, -32'd1478},
{-32'd149, 32'd4484, 32'd8941, -32'd5640},
{32'd4153, -32'd2668, -32'd4209, 32'd1073},
{-32'd4279, -32'd3272, -32'd6986, 32'd3488},
{-32'd15742, -32'd3738, 32'd9574, -32'd5572},
{-32'd4810, -32'd1682, -32'd12524, -32'd4014},
{-32'd2474, 32'd718, -32'd6859, 32'd548},
{32'd3605, -32'd5343, 32'd3632, -32'd3494},
{-32'd4543, 32'd6159, 32'd3663, 32'd1577},
{32'd130, 32'd1535, -32'd1341, 32'd5227},
{32'd770, 32'd8176, -32'd7228, 32'd7131},
{-32'd2700, -32'd3552, 32'd2259, 32'd7056},
{32'd1439, 32'd77, -32'd1860, -32'd3304},
{32'd6231, -32'd2418, 32'd72, -32'd3492},
{32'd16775, -32'd6579, -32'd10992, 32'd2933},
{32'd741, 32'd3248, -32'd7162, -32'd3832},
{32'd2088, 32'd2860, 32'd8472, -32'd3261},
{32'd14227, 32'd5883, 32'd5346, 32'd4891},
{32'd2880, -32'd719, 32'd7416, -32'd869},
{-32'd7703, 32'd4403, -32'd44, -32'd5291},
{32'd12399, 32'd1163, -32'd3423, -32'd2442},
{-32'd14144, 32'd4745, -32'd440, -32'd592},
{32'd1764, -32'd7993, -32'd3819, -32'd2191},
{32'd6199, -32'd7931, -32'd7451, 32'd3297},
{-32'd6280, -32'd4336, -32'd4115, 32'd1074},
{32'd6024, 32'd10417, 32'd19872, 32'd3558},
{-32'd7426, -32'd10254, 32'd2701, -32'd434},
{32'd7922, -32'd812, -32'd9225, 32'd235},
{32'd13373, 32'd10916, 32'd9569, 32'd1199},
{-32'd8024, 32'd358, 32'd386, 32'd5318},
{32'd3084, -32'd8941, -32'd3272, 32'd5132},
{-32'd8811, 32'd6116, -32'd7909, 32'd6156},
{-32'd7801, 32'd4417, 32'd4063, 32'd12883},
{32'd4635, -32'd5789, -32'd235, -32'd4705},
{-32'd2141, 32'd808, 32'd2358, 32'd2202},
{32'd595, 32'd3835, -32'd4711, -32'd6767},
{32'd1185, 32'd5843, -32'd922, 32'd3003},
{-32'd6044, -32'd7561, 32'd5136, 32'd7921},
{-32'd4238, 32'd9010, -32'd1880, -32'd7923},
{-32'd6680, -32'd1839, 32'd4231, -32'd16},
{-32'd1144, -32'd7968, 32'd856, -32'd240},
{32'd2123, -32'd6073, 32'd829, -32'd2262},
{-32'd4087, -32'd1943, -32'd9931, -32'd3347},
{32'd1839, -32'd995, -32'd2146, -32'd2789},
{32'd184, 32'd7771, 32'd1406, 32'd2784},
{32'd432, -32'd5327, -32'd3676, 32'd771},
{32'd19804, -32'd3034, -32'd2853, -32'd4039},
{32'd558, -32'd5773, 32'd9185, -32'd3387},
{32'd2793, -32'd3143, 32'd5847, 32'd220},
{-32'd1949, -32'd6539, -32'd7369, -32'd7646},
{32'd3939, 32'd1792, -32'd445, 32'd3994},
{-32'd830, -32'd6927, 32'd595, 32'd1440},
{32'd3164, -32'd10253, -32'd4742, -32'd16554},
{-32'd5536, -32'd3709, -32'd2853, 32'd8197},
{-32'd12844, 32'd409, -32'd20700, -32'd9115},
{32'd1301, 32'd2334, -32'd5963, -32'd520},
{-32'd5187, 32'd3337, -32'd383, 32'd705},
{32'd5400, -32'd2268, -32'd4190, -32'd4086},
{32'd9663, 32'd2892, -32'd3757, 32'd5134},
{-32'd3094, -32'd274, -32'd25, -32'd4122},
{32'd9277, -32'd466, -32'd333, 32'd7141},
{-32'd4963, -32'd3943, 32'd3486, -32'd4663},
{-32'd346, -32'd3904, -32'd7496, 32'd1149},
{-32'd9237, -32'd13539, -32'd971, -32'd456},
{-32'd3233, -32'd4449, -32'd3356, 32'd3827},
{32'd4293, 32'd10355, 32'd6491, 32'd4580},
{32'd690, 32'd83, 32'd4092, -32'd10067},
{32'd9244, -32'd466, -32'd4146, -32'd8572},
{32'd8129, -32'd12649, -32'd13583, 32'd239},
{32'd4280, -32'd10283, 32'd183, -32'd13615},
{32'd13225, -32'd3889, 32'd161, 32'd1741},
{32'd7476, 32'd3531, 32'd1869, 32'd1610},
{-32'd7586, -32'd12179, -32'd790, 32'd1273},
{32'd8896, -32'd6635, -32'd7820, -32'd12103},
{32'd567, -32'd6290, 32'd5291, 32'd9635},
{32'd5445, 32'd2404, 32'd1835, 32'd13271},
{-32'd11984, -32'd4309, 32'd3807, -32'd12469},
{-32'd7216, 32'd2413, -32'd3896, 32'd15225},
{-32'd3615, -32'd7696, 32'd2263, -32'd7027},
{32'd10953, -32'd2938, 32'd563, 32'd3861},
{32'd21674, -32'd28, 32'd3583, -32'd920},
{-32'd443, 32'd13677, 32'd3808, 32'd1548},
{-32'd7411, -32'd7661, 32'd459, -32'd8966},
{-32'd700, -32'd1240, 32'd7966, -32'd3883},
{-32'd3300, -32'd21, -32'd8638, 32'd5749},
{32'd7994, -32'd8168, -32'd13861, 32'd1351},
{-32'd601, 32'd2544, -32'd4483, -32'd2669},
{32'd3568, -32'd7605, -32'd5390, 32'd5845},
{32'd6582, -32'd3702, -32'd7593, 32'd3624},
{32'd749, 32'd3296, -32'd12152, -32'd2514},
{32'd5595, -32'd4805, 32'd12613, -32'd641},
{-32'd4182, 32'd9096, -32'd3969, -32'd3186},
{-32'd8117, -32'd572, 32'd139, 32'd266},
{-32'd3644, 32'd6031, -32'd2921, 32'd7722},
{32'd905, 32'd6065, -32'd13951, -32'd1617},
{32'd2111, -32'd510, -32'd977, -32'd5757},
{32'd944, -32'd3241, -32'd1403, -32'd3711},
{-32'd9591, -32'd8935, -32'd267, 32'd15101},
{-32'd801, 32'd5121, 32'd3501, -32'd9457},
{32'd955, -32'd144, -32'd830, 32'd5075},
{32'd381, 32'd5747, -32'd6258, 32'd1895},
{32'd5592, 32'd2266, 32'd14240, 32'd9585},
{-32'd5376, -32'd3824, -32'd6751, -32'd4198},
{32'd663, -32'd1571, 32'd5225, 32'd119},
{32'd17170, -32'd176, -32'd10649, -32'd1020},
{-32'd4701, 32'd4489, 32'd5190, 32'd515},
{-32'd10586, -32'd451, 32'd7160, -32'd6485},
{-32'd11711, 32'd2897, 32'd4528, 32'd356},
{-32'd5933, -32'd9725, 32'd8684, 32'd4349},
{32'd8427, -32'd2287, -32'd5566, -32'd4505},
{32'd4039, 32'd9478, 32'd1257, -32'd4354},
{-32'd4128, -32'd2959, 32'd4807, -32'd5986},
{-32'd69, 32'd11855, -32'd1024, -32'd11139},
{-32'd2248, 32'd4389, 32'd2480, 32'd691},
{-32'd5963, -32'd15247, -32'd3338, -32'd5974},
{32'd93, -32'd2987, 32'd9543, -32'd7379},
{32'd5481, 32'd10779, 32'd4607, 32'd2028},
{-32'd4631, -32'd2647, 32'd6611, -32'd4537},
{-32'd6149, -32'd7485, -32'd8267, -32'd5713},
{-32'd903, 32'd5372, 32'd10369, -32'd513},
{-32'd3051, 32'd5419, -32'd15278, -32'd4479},
{-32'd3161, 32'd10855, 32'd10344, -32'd1335},
{-32'd2348, -32'd6082, 32'd4265, -32'd3132},
{-32'd2102, 32'd3319, -32'd324, 32'd1222},
{32'd562, -32'd2439, 32'd10941, -32'd13609},
{32'd1336, -32'd12003, 32'd1422, 32'd4440},
{32'd432, -32'd12910, -32'd3654, -32'd4864},
{-32'd3198, -32'd1509, 32'd1000, -32'd5990},
{32'd5573, -32'd2770, 32'd6834, -32'd12456},
{32'd9744, 32'd4402, 32'd10738, -32'd3356},
{-32'd10465, -32'd8215, 32'd1417, -32'd4451},
{32'd4527, -32'd6067, 32'd3804, 32'd1323},
{32'd4392, -32'd6074, 32'd3513, -32'd7960},
{-32'd5990, 32'd9286, -32'd2729, -32'd518},
{-32'd4405, -32'd7793, -32'd5906, 32'd3337},
{-32'd1848, -32'd4766, 32'd2093, -32'd9727},
{32'd4477, -32'd7500, -32'd593, -32'd3500},
{-32'd8891, 32'd4628, -32'd12962, -32'd1138},
{32'd8703, 32'd6401, 32'd8629, 32'd6368},
{32'd13301, -32'd5255, 32'd2605, 32'd1468},
{-32'd3379, -32'd2125, 32'd2793, 32'd6542},
{-32'd3945, -32'd7826, -32'd1547, 32'd12006},
{-32'd724, 32'd5366, -32'd5053, 32'd2452},
{-32'd4269, 32'd7028, 32'd3428, 32'd3183},
{-32'd11430, -32'd7050, -32'd13111, -32'd1471},
{32'd952, -32'd10857, -32'd1080, -32'd1841},
{32'd721, -32'd1027, -32'd673, 32'd2502},
{-32'd4922, -32'd3, 32'd1113, 32'd5457},
{32'd6816, 32'd7880, 32'd3823, 32'd3581},
{32'd7200, -32'd2848, -32'd1579, -32'd12318},
{-32'd4500, 32'd2331, -32'd1295, -32'd1836},
{-32'd6324, 32'd3805, 32'd2902, -32'd2302},
{-32'd1031, 32'd14557, -32'd3154, 32'd3982},
{32'd3966, 32'd10473, 32'd701, -32'd9491},
{32'd3895, -32'd321, 32'd1478, -32'd1331},
{32'd7686, -32'd7832, -32'd8160, -32'd2905},
{32'd5824, -32'd177, 32'd3634, 32'd10200},
{-32'd6623, -32'd13034, -32'd2354, -32'd4460},
{32'd828, -32'd8836, -32'd3813, 32'd1388},
{-32'd9623, 32'd2388, -32'd5281, -32'd10509},
{32'd3749, -32'd7751, 32'd4258, 32'd5222},
{-32'd11286, -32'd4831, -32'd1170, 32'd4468},
{-32'd5047, 32'd3542, -32'd2218, -32'd2938},
{32'd12981, 32'd3612, 32'd9397, 32'd8036},
{32'd5671, -32'd5877, -32'd10061, 32'd255},
{32'd921, -32'd2918, 32'd1999, -32'd4859},
{32'd7105, -32'd644, -32'd2039, -32'd8832},
{-32'd3619, -32'd4273, -32'd710, 32'd3914},
{-32'd3932, 32'd2246, -32'd862, 32'd3019},
{32'd6757, 32'd1526, 32'd3881, -32'd25},
{-32'd1218, -32'd1113, -32'd3080, 32'd2036},
{-32'd54, -32'd13344, -32'd6700, -32'd4026}
},
{{32'd2982, 32'd13656, 32'd4765, 32'd6099},
{-32'd10520, -32'd5936, -32'd8741, -32'd2853},
{32'd5133, -32'd821, 32'd13319, -32'd8579},
{32'd245, 32'd4289, -32'd6493, 32'd8301},
{32'd14490, 32'd3675, 32'd8428, -32'd2870},
{-32'd7730, 32'd5448, -32'd7210, 32'd2125},
{32'd9475, -32'd10379, 32'd18033, -32'd16592},
{32'd4726, 32'd7725, -32'd6492, -32'd10288},
{32'd9231, -32'd4175, -32'd5808, 32'd1479},
{32'd7598, 32'd5270, 32'd7489, 32'd13987},
{-32'd6480, -32'd9220, 32'd14065, -32'd3113},
{32'd9685, -32'd4605, -32'd5145, -32'd4888},
{32'd10099, -32'd7410, -32'd6261, 32'd9255},
{-32'd2681, 32'd2338, 32'd10775, -32'd612},
{-32'd6146, -32'd597, -32'd3466, -32'd1889},
{-32'd1096, -32'd1913, 32'd1591, -32'd7470},
{32'd4897, 32'd4355, 32'd1629, -32'd641},
{32'd970, 32'd23495, 32'd4539, 32'd6760},
{32'd1023, -32'd3715, 32'd5915, -32'd8571},
{32'd14985, 32'd4913, 32'd3486, 32'd1773},
{32'd9969, -32'd11328, -32'd2199, 32'd4365},
{-32'd3861, 32'd4675, 32'd2111, 32'd536},
{-32'd3475, -32'd10425, -32'd11347, -32'd1948},
{-32'd2892, 32'd5093, 32'd3609, -32'd5103},
{32'd1515, -32'd2106, 32'd5016, 32'd5770},
{32'd14895, 32'd853, 32'd5597, -32'd10649},
{-32'd8988, -32'd1701, -32'd6111, -32'd7903},
{32'd3186, -32'd3478, -32'd878, -32'd9550},
{32'd2980, 32'd3149, 32'd10944, 32'd2763},
{32'd440, 32'd613, 32'd9001, 32'd4426},
{32'd8431, 32'd12315, 32'd6133, -32'd5566},
{-32'd9643, 32'd7766, 32'd1556, -32'd5747},
{32'd7354, -32'd8399, 32'd12457, -32'd434},
{32'd5110, 32'd1301, 32'd11078, -32'd9724},
{32'd6432, 32'd18784, -32'd285, 32'd11277},
{-32'd5967, 32'd17719, 32'd2371, -32'd1969},
{-32'd4600, 32'd2420, 32'd852, -32'd22701},
{-32'd5235, 32'd8564, 32'd3440, 32'd6105},
{32'd5707, -32'd7943, 32'd4677, 32'd5764},
{-32'd22060, -32'd9867, -32'd10866, 32'd480},
{-32'd753, -32'd9837, 32'd2744, -32'd7281},
{32'd1450, 32'd9072, -32'd597, -32'd5826},
{32'd333, 32'd10816, -32'd845, 32'd10091},
{-32'd5999, -32'd9675, -32'd6834, -32'd12485},
{-32'd3826, 32'd3785, -32'd5549, 32'd2930},
{-32'd10784, -32'd3281, -32'd4843, -32'd5351},
{32'd3737, 32'd10248, 32'd5203, 32'd4193},
{32'd2517, 32'd2575, 32'd769, -32'd5473},
{32'd14831, -32'd367, 32'd6593, 32'd848},
{-32'd6693, 32'd10086, -32'd10005, 32'd10030},
{32'd5693, -32'd6638, -32'd1864, -32'd1204},
{-32'd7113, 32'd3478, -32'd6697, -32'd823},
{32'd4986, 32'd3050, 32'd1728, -32'd1624},
{-32'd1474, 32'd8086, -32'd4347, -32'd666},
{32'd12436, 32'd2700, -32'd6006, -32'd2958},
{-32'd11333, -32'd13853, -32'd2224, 32'd2171},
{-32'd5704, -32'd8031, -32'd2267, 32'd3920},
{32'd3942, -32'd4524, -32'd5674, -32'd6626},
{-32'd11592, 32'd4259, -32'd5900, 32'd2932},
{-32'd10866, 32'd713, -32'd7265, 32'd5627},
{32'd6564, 32'd6045, -32'd1036, -32'd3439},
{-32'd899, -32'd2636, 32'd6254, -32'd3461},
{-32'd7362, -32'd4183, 32'd1420, -32'd5176},
{32'd6247, -32'd1511, -32'd5226, 32'd7898},
{-32'd169, 32'd5399, 32'd575, 32'd8854},
{32'd11507, 32'd5659, -32'd4904, 32'd5612},
{-32'd123, -32'd10009, -32'd351, -32'd2331},
{-32'd1571, 32'd6891, -32'd10814, -32'd4255},
{32'd284, 32'd833, 32'd3576, 32'd683},
{-32'd122, 32'd12293, -32'd11084, -32'd9553},
{-32'd14367, -32'd1383, -32'd1632, -32'd5150},
{-32'd11621, 32'd10532, 32'd1017, -32'd3004},
{-32'd20848, -32'd2317, 32'd4799, -32'd8313},
{32'd5938, -32'd20243, -32'd4965, 32'd9738},
{32'd12346, 32'd3476, 32'd6074, 32'd7725},
{-32'd4713, 32'd11108, -32'd2394, -32'd10362},
{32'd2075, 32'd6018, -32'd6233, 32'd276},
{32'd603, -32'd3410, 32'd4780, -32'd2152},
{32'd4774, 32'd10788, 32'd3607, -32'd5992},
{-32'd3088, -32'd6681, -32'd7847, -32'd6641},
{32'd1535, 32'd5776, 32'd293, -32'd6815},
{-32'd8414, 32'd527, -32'd8255, -32'd985},
{-32'd11423, -32'd17563, -32'd5233, -32'd7928},
{-32'd10343, 32'd3046, 32'd2379, -32'd4763},
{-32'd1710, -32'd5832, 32'd4980, 32'd6761},
{32'd3714, -32'd4850, 32'd3609, 32'd5566},
{32'd1726, 32'd14138, 32'd5547, -32'd3364},
{-32'd2892, -32'd9877, 32'd8761, 32'd1740},
{32'd9144, 32'd7142, 32'd2354, -32'd14553},
{-32'd3806, 32'd2281, 32'd220, 32'd651},
{32'd863, -32'd6383, 32'd3330, 32'd6123},
{-32'd8660, -32'd16499, -32'd6712, -32'd628},
{32'd4774, 32'd13362, 32'd310, 32'd9399},
{32'd8367, 32'd8936, 32'd7321, 32'd15667},
{32'd5949, 32'd9838, -32'd5799, 32'd2131},
{-32'd12683, 32'd1172, 32'd6307, 32'd10112},
{32'd10706, 32'd10003, 32'd8305, 32'd4849},
{32'd3821, 32'd12698, 32'd4017, -32'd623},
{-32'd115, -32'd6381, 32'd13742, -32'd8184},
{32'd2161, 32'd17941, 32'd9118, 32'd12354},
{-32'd3033, -32'd16146, -32'd3052, 32'd11131},
{-32'd10761, 32'd12379, -32'd12768, -32'd7122},
{-32'd2649, -32'd13400, -32'd9337, -32'd5404},
{-32'd3918, 32'd17904, -32'd2889, 32'd5726},
{32'd13973, 32'd6861, -32'd5779, 32'd5195},
{32'd1142, -32'd4853, -32'd3458, 32'd205},
{-32'd8998, 32'd2202, -32'd10135, -32'd3823},
{32'd3381, 32'd3958, 32'd1686, 32'd12387},
{32'd165, 32'd8318, -32'd3234, 32'd4009},
{32'd202, 32'd6704, -32'd6603, -32'd4780},
{-32'd12465, 32'd2526, 32'd1611, -32'd17371},
{-32'd8885, -32'd5764, 32'd13791, 32'd2957},
{-32'd1776, 32'd9168, 32'd3152, 32'd1357},
{32'd763, 32'd5261, 32'd8475, -32'd13274},
{-32'd2490, 32'd4097, -32'd16075, -32'd1876},
{-32'd7788, -32'd8675, -32'd13462, 32'd1498},
{32'd9746, 32'd4996, -32'd2456, -32'd795},
{-32'd14154, 32'd1761, 32'd9150, 32'd2999},
{-32'd15620, 32'd7924, -32'd7931, 32'd6680},
{32'd6529, 32'd3661, 32'd2354, 32'd9436},
{32'd16521, -32'd1548, -32'd1498, -32'd2554},
{32'd499, 32'd458, 32'd8547, -32'd12522},
{32'd18800, 32'd1942, -32'd3093, 32'd3399},
{-32'd4186, 32'd190, 32'd3445, -32'd2281},
{32'd6014, 32'd2106, 32'd112, -32'd2942},
{-32'd11991, 32'd12983, 32'd3116, 32'd1482},
{-32'd7916, 32'd11399, -32'd13116, -32'd5360},
{-32'd4374, -32'd304, -32'd9737, -32'd1275},
{-32'd16291, -32'd5987, -32'd2116, -32'd1328},
{32'd9415, -32'd9658, 32'd6940, -32'd11776},
{-32'd2197, 32'd19144, 32'd1738, 32'd3836},
{-32'd12062, -32'd2384, -32'd9680, -32'd5079},
{32'd2087, -32'd6296, -32'd3857, -32'd4345},
{-32'd3400, -32'd4128, -32'd4983, 32'd5932},
{32'd4468, 32'd6092, -32'd7448, -32'd10596},
{-32'd11312, -32'd13826, 32'd7553, -32'd1344},
{32'd4926, -32'd894, -32'd5608, -32'd11780},
{32'd699, 32'd1929, -32'd5227, 32'd5753},
{32'd8751, -32'd8990, 32'd11462, -32'd5733},
{32'd1765, -32'd11110, -32'd7203, -32'd5900},
{-32'd5473, -32'd4050, -32'd7327, 32'd9392},
{-32'd3944, -32'd10242, -32'd6970, -32'd5550},
{-32'd456, 32'd9515, 32'd9914, -32'd1812},
{-32'd6822, -32'd9151, 32'd8688, 32'd395},
{32'd2596, 32'd7449, 32'd9554, 32'd11591},
{-32'd6324, -32'd6985, -32'd3346, 32'd917},
{-32'd8411, 32'd5310, 32'd2950, 32'd2152},
{-32'd1106, -32'd1958, 32'd4756, -32'd2393},
{-32'd4618, -32'd10087, -32'd7869, 32'd1723},
{-32'd3122, -32'd762, -32'd4279, -32'd8369},
{-32'd2627, -32'd139, 32'd3036, -32'd24674},
{-32'd5237, 32'd1707, 32'd13600, 32'd11386},
{-32'd434, -32'd6128, -32'd420, -32'd1896},
{32'd1518, 32'd14408, -32'd3644, -32'd6877},
{-32'd16496, -32'd7496, -32'd4625, -32'd8553},
{32'd5048, -32'd11242, -32'd8393, -32'd14818},
{32'd7230, -32'd7992, -32'd10670, 32'd913},
{32'd5544, -32'd398, -32'd818, -32'd5389},
{-32'd5586, 32'd3295, -32'd349, 32'd6518},
{32'd3038, 32'd5469, 32'd9289, 32'd7691},
{-32'd7190, 32'd21343, -32'd3516, 32'd3307},
{32'd1324, -32'd1734, -32'd1956, -32'd3413},
{-32'd8548, 32'd15377, -32'd2361, 32'd9844},
{32'd6185, 32'd14321, 32'd7270, 32'd9034},
{-32'd1642, -32'd1935, -32'd3735, 32'd2366},
{-32'd17765, -32'd7756, 32'd4626, 32'd8779},
{32'd10008, -32'd6669, -32'd3644, 32'd4115},
{-32'd4291, 32'd16224, -32'd2094, -32'd3160},
{32'd3929, 32'd12592, 32'd5259, 32'd659},
{32'd8870, -32'd11558, 32'd3187, -32'd10301},
{-32'd7759, -32'd2506, -32'd235, 32'd6593},
{-32'd9360, -32'd18079, -32'd2438, -32'd1645},
{32'd4883, 32'd5081, -32'd895, 32'd14645},
{32'd805, 32'd3259, 32'd1252, -32'd6564},
{32'd8309, 32'd17450, 32'd1714, 32'd6209},
{-32'd2168, -32'd7883, 32'd12818, 32'd5268},
{32'd5316, -32'd8262, 32'd73, -32'd8658},
{-32'd10255, -32'd10452, 32'd4357, 32'd284},
{32'd5527, 32'd10653, -32'd4879, 32'd3495},
{-32'd9573, -32'd5877, -32'd4916, -32'd14489},
{-32'd5442, -32'd6258, -32'd6708, 32'd3831},
{-32'd6220, 32'd5061, -32'd8504, -32'd6810},
{-32'd2647, -32'd9217, 32'd7334, 32'd4305},
{-32'd11016, 32'd16635, -32'd10229, 32'd1215},
{32'd4980, -32'd5261, 32'd1156, 32'd8202},
{32'd4521, -32'd12527, 32'd1946, -32'd1438},
{-32'd6628, 32'd2825, -32'd5766, 32'd12941},
{-32'd17934, 32'd2116, -32'd12632, 32'd23803},
{-32'd988, -32'd7790, 32'd883, 32'd11065},
{-32'd9920, -32'd1492, -32'd2779, -32'd7291},
{-32'd4830, 32'd6311, -32'd4369, -32'd2924},
{32'd461, -32'd5193, -32'd5062, -32'd1515},
{-32'd8917, 32'd6822, -32'd11772, 32'd7701},
{32'd6042, 32'd4586, -32'd12938, -32'd5068},
{-32'd4079, -32'd2989, 32'd2901, -32'd2743},
{-32'd840, 32'd7568, -32'd6, -32'd6890},
{-32'd20735, 32'd6745, 32'd323, -32'd7452},
{-32'd1302, -32'd9560, 32'd5649, 32'd7184},
{32'd3567, -32'd10057, 32'd3326, -32'd5047},
{-32'd3846, 32'd2565, 32'd4319, -32'd261},
{-32'd10388, -32'd2414, -32'd4108, -32'd8377},
{-32'd7741, 32'd3860, -32'd5757, -32'd3062},
{32'd15061, -32'd8742, 32'd7180, -32'd10360},
{-32'd1239, 32'd2872, -32'd151, 32'd8422},
{-32'd1171, 32'd4142, -32'd887, -32'd2021},
{-32'd1861, 32'd8842, 32'd427, -32'd1924},
{-32'd7795, -32'd3195, 32'd2449, 32'd9023},
{32'd1771, 32'd6770, 32'd3956, -32'd5131},
{32'd9688, -32'd816, 32'd8955, -32'd12129},
{32'd17405, 32'd26593, 32'd6803, -32'd2167},
{-32'd8393, -32'd4806, -32'd4469, -32'd3131},
{32'd3104, 32'd5516, 32'd6316, 32'd4060},
{32'd2662, 32'd605, -32'd3729, -32'd5248},
{-32'd4316, 32'd516, 32'd6370, -32'd741},
{-32'd7647, -32'd10574, -32'd538, 32'd4979},
{32'd7513, -32'd5554, -32'd6402, 32'd4355},
{-32'd14666, 32'd5909, -32'd11373, -32'd3928},
{32'd5933, -32'd7743, -32'd261, -32'd1749},
{-32'd2479, 32'd6025, -32'd2795, 32'd13828},
{32'd2352, 32'd4647, -32'd9685, 32'd3600},
{-32'd16879, -32'd884, -32'd5046, 32'd908},
{32'd4633, 32'd1383, -32'd4984, -32'd1049},
{32'd2319, 32'd12433, -32'd240, -32'd8288},
{32'd2743, -32'd17002, 32'd5759, 32'd1113},
{32'd6667, -32'd5547, 32'd5991, -32'd5312},
{-32'd9117, -32'd4528, -32'd3637, -32'd2117},
{-32'd14337, 32'd9090, 32'd314, -32'd4631},
{32'd2309, -32'd5478, -32'd7782, -32'd4221},
{32'd5506, -32'd2878, -32'd2905, -32'd4500},
{32'd6645, 32'd5382, -32'd1746, -32'd7314},
{-32'd13730, -32'd1954, 32'd746, -32'd5066},
{-32'd10217, -32'd2111, -32'd2936, -32'd8036},
{32'd2308, -32'd15908, 32'd10276, -32'd7021},
{-32'd4995, 32'd11029, -32'd8161, 32'd5016},
{-32'd9158, -32'd2712, 32'd2139, 32'd911},
{-32'd12230, 32'd3927, 32'd4036, -32'd2555},
{-32'd11128, -32'd12829, 32'd16415, 32'd2689},
{-32'd3402, -32'd6816, 32'd6582, -32'd1497},
{32'd1974, 32'd3404, -32'd2621, -32'd6008},
{32'd9231, 32'd5732, -32'd2125, -32'd8543},
{-32'd912, -32'd7719, -32'd7241, 32'd529},
{32'd2703, 32'd1889, -32'd861, -32'd2687},
{-32'd3350, 32'd821, -32'd4283, -32'd14604},
{-32'd7692, -32'd15335, -32'd3909, -32'd1176},
{32'd2849, 32'd3347, 32'd5499, 32'd5613},
{32'd4112, 32'd17970, 32'd7359, -32'd1215},
{-32'd10614, -32'd8356, 32'd1455, -32'd1317},
{-32'd10262, 32'd12140, 32'd2134, 32'd11306},
{32'd3065, 32'd9237, 32'd865, 32'd1641},
{-32'd4940, -32'd1469, -32'd5860, -32'd1423},
{-32'd3023, 32'd2144, 32'd3777, -32'd2449},
{32'd3514, 32'd4223, -32'd2034, 32'd7452},
{-32'd2081, 32'd2647, 32'd943, 32'd5949},
{-32'd223, -32'd1849, -32'd7896, 32'd10018},
{-32'd5311, -32'd1624, 32'd1183, 32'd1969},
{32'd4361, 32'd2048, -32'd3222, 32'd7174},
{32'd3923, -32'd4728, -32'd1748, 32'd7165},
{32'd8186, 32'd768, -32'd7375, 32'd15123},
{-32'd1160, -32'd10489, 32'd1446, 32'd2668},
{-32'd2401, 32'd6592, 32'd5921, -32'd10227},
{-32'd992, -32'd3496, -32'd1618, 32'd7736},
{-32'd5707, 32'd15122, 32'd3412, 32'd5643},
{-32'd4616, 32'd8564, 32'd7177, -32'd9410},
{-32'd2973, -32'd4091, -32'd995, -32'd10421},
{32'd4298, -32'd983, 32'd259, -32'd4708},
{-32'd5491, -32'd22164, 32'd3584, 32'd3002},
{32'd3456, 32'd2623, -32'd7123, 32'd2448},
{32'd939, 32'd6817, 32'd2416, -32'd6735},
{-32'd1758, 32'd1118, 32'd6613, -32'd11191},
{-32'd8620, 32'd10560, 32'd6323, 32'd5678},
{-32'd2212, -32'd5259, 32'd2192, 32'd6208},
{32'd5020, -32'd5042, -32'd3802, -32'd5642},
{32'd3278, 32'd14959, 32'd7875, -32'd3578},
{-32'd7110, -32'd4794, -32'd13432, 32'd3572},
{-32'd5332, 32'd2241, 32'd2991, 32'd6215},
{-32'd7517, -32'd9291, 32'd2943, -32'd15586},
{32'd11295, 32'd5675, 32'd4209, 32'd15970},
{-32'd8205, 32'd1599, 32'd421, -32'd7206},
{-32'd33, -32'd8043, 32'd3216, -32'd12556},
{-32'd2303, 32'd1743, -32'd2377, -32'd1951},
{32'd9741, 32'd578, -32'd4661, 32'd1968},
{-32'd3929, -32'd719, -32'd3212, 32'd10137},
{32'd7218, -32'd10171, 32'd7294, -32'd4968},
{32'd4411, -32'd7795, -32'd5799, 32'd6245},
{32'd5623, -32'd2425, -32'd2514, 32'd985},
{-32'd5412, -32'd10720, -32'd2579, -32'd4103},
{32'd2264, 32'd5720, 32'd2226, 32'd5352},
{-32'd5510, 32'd2175, 32'd2021, 32'd1216},
{-32'd536, 32'd4857, 32'd1615, 32'd4161},
{-32'd5806, 32'd11560, 32'd3307, -32'd7163},
{32'd8999, 32'd3143, -32'd7036, -32'd11828},
{32'd8202, 32'd2733, 32'd2516, 32'd8697},
{-32'd12429, -32'd8579, -32'd2680, 32'd28},
{32'd504, -32'd1274, 32'd12100, -32'd5445},
{32'd5024, -32'd14924, 32'd3008, -32'd3436},
{-32'd1643, -32'd1249, -32'd1597, -32'd6148},
{-32'd9468, -32'd3245, -32'd7187, 32'd2710},
{32'd7051, 32'd10326, 32'd4338, 32'd12471},
{32'd6641, -32'd3839, 32'd362, 32'd3293},
{32'd1130, -32'd6553, 32'd8837, -32'd4235}
},
{{32'd12292, 32'd8566, 32'd3651, 32'd2320},
{-32'd11076, -32'd5187, 32'd312, -32'd3881},
{32'd3103, 32'd1689, 32'd7751, 32'd3996},
{-32'd14094, 32'd5573, 32'd4388, 32'd9042},
{-32'd5629, -32'd1944, 32'd2836, -32'd495},
{32'd5568, -32'd6284, 32'd11098, 32'd438},
{32'd866, 32'd6969, -32'd2437, 32'd3559},
{32'd1136, -32'd637, 32'd10795, -32'd190},
{-32'd968, 32'd3409, -32'd126, 32'd1440},
{32'd3095, 32'd10240, 32'd2287, 32'd5458},
{-32'd6911, 32'd312, 32'd6678, 32'd2153},
{-32'd2600, 32'd549, -32'd871, -32'd7471},
{-32'd2264, 32'd772, -32'd9263, 32'd1549},
{-32'd11504, 32'd192, 32'd1331, -32'd2715},
{-32'd6215, -32'd170, -32'd2959, 32'd297},
{32'd1840, -32'd11621, -32'd7452, -32'd7155},
{32'd4604, -32'd534, 32'd10270, 32'd6041},
{-32'd823, 32'd8018, -32'd201, 32'd6535},
{-32'd10136, 32'd1818, 32'd8191, 32'd5734},
{32'd3809, -32'd4352, 32'd6564, 32'd4606},
{-32'd10584, 32'd1717, 32'd7356, 32'd5919},
{-32'd679, -32'd4314, 32'd341, 32'd1370},
{32'd8352, -32'd9064, -32'd2610, -32'd3200},
{-32'd5378, -32'd2977, -32'd4869, -32'd6433},
{-32'd437, 32'd5336, -32'd1796, -32'd14},
{-32'd3505, 32'd4172, 32'd13882, 32'd7196},
{-32'd930, 32'd4702, 32'd13036, -32'd2374},
{32'd2588, -32'd3459, -32'd922, 32'd89},
{32'd2143, 32'd1033, 32'd10404, 32'd1518},
{32'd16855, 32'd6026, -32'd14913, -32'd5259},
{-32'd1188, 32'd1413, 32'd2375, 32'd4311},
{32'd2672, -32'd10257, 32'd3930, -32'd4377},
{32'd7588, -32'd801, -32'd1733, 32'd4275},
{32'd3933, -32'd170, -32'd12593, -32'd5300},
{32'd10890, 32'd7594, 32'd4938, 32'd3174},
{32'd5047, -32'd4380, -32'd8881, 32'd7910},
{32'd6874, -32'd1320, 32'd5195, -32'd1512},
{-32'd7745, 32'd2363, -32'd5344, -32'd603},
{32'd6367, -32'd1609, -32'd11556, -32'd388},
{32'd1393, 32'd1091, 32'd2260, 32'd2533},
{32'd3781, 32'd2461, -32'd6082, -32'd7571},
{32'd3500, 32'd4372, -32'd3664, 32'd5193},
{-32'd1054, 32'd1733, -32'd3978, 32'd3133},
{-32'd7223, -32'd6670, -32'd10557, -32'd8015},
{32'd3665, 32'd1703, -32'd10378, -32'd3638},
{-32'd609, -32'd3913, -32'd16692, -32'd8525},
{32'd7478, -32'd7198, 32'd1816, -32'd1059},
{-32'd1350, -32'd5019, -32'd3030, -32'd2974},
{32'd5653, 32'd76, 32'd1180, 32'd5506},
{32'd9318, -32'd10860, -32'd3824, -32'd6288},
{-32'd6775, 32'd1559, -32'd98, 32'd1428},
{32'd5035, -32'd3403, -32'd12695, -32'd5140},
{-32'd2533, -32'd419, 32'd6961, 32'd2134},
{-32'd13510, 32'd1670, -32'd4129, 32'd309},
{32'd2022, 32'd7442, -32'd2701, -32'd4873},
{32'd3989, -32'd4533, -32'd3322, -32'd1498},
{32'd3764, 32'd753, 32'd1834, 32'd8293},
{32'd3205, -32'd5448, 32'd1741, 32'd1495},
{-32'd5077, -32'd5751, 32'd2841, -32'd4007},
{32'd11046, 32'd926, 32'd322, -32'd1487},
{-32'd9178, -32'd2606, -32'd614, 32'd5522},
{32'd579, -32'd6766, 32'd6703, -32'd898},
{-32'd6919, -32'd2034, 32'd2972, 32'd1504},
{32'd9553, 32'd569, 32'd3382, 32'd2569},
{32'd4100, -32'd2980, -32'd13078, -32'd7745},
{-32'd5886, 32'd11334, -32'd585, 32'd5707},
{-32'd4958, -32'd4342, 32'd4792, -32'd6676},
{32'd963, -32'd2287, -32'd1614, -32'd4493},
{32'd6769, -32'd537, -32'd5405, -32'd2567},
{-32'd2064, -32'd5490, 32'd4940, -32'd2940},
{32'd6818, 32'd2057, -32'd5743, -32'd8434},
{32'd2239, 32'd572, -32'd4183, -32'd1034},
{-32'd5013, 32'd592, -32'd5964, -32'd7942},
{32'd5624, -32'd5367, -32'd3029, 32'd3855},
{32'd9574, 32'd10034, -32'd2308, -32'd785},
{32'd7544, 32'd5534, -32'd3094, -32'd6379},
{-32'd7819, -32'd3433, -32'd1701, -32'd3921},
{-32'd188, -32'd6669, 32'd10691, 32'd2520},
{-32'd815, 32'd4061, -32'd10318, 32'd3635},
{-32'd7792, 32'd8763, 32'd6193, 32'd5226},
{32'd2289, -32'd1141, -32'd1718, -32'd1086},
{-32'd7140, -32'd8173, -32'd6271, 32'd1724},
{-32'd3910, -32'd5648, 32'd5133, 32'd4562},
{-32'd3564, 32'd10239, -32'd15421, -32'd9839},
{-32'd6806, 32'd5706, -32'd13803, -32'd5109},
{32'd8295, -32'd2934, -32'd3667, -32'd6484},
{32'd11597, -32'd2078, -32'd6104, 32'd1560},
{-32'd3109, -32'd7819, -32'd428, -32'd2453},
{32'd802, -32'd1928, -32'd1269, -32'd13},
{32'd3501, 32'd1506, 32'd682, -32'd7111},
{32'd852, 32'd5808, -32'd7473, 32'd1727},
{-32'd6311, -32'd3578, -32'd14113, 32'd4026},
{-32'd826, -32'd1553, 32'd494, 32'd3397},
{32'd8156, -32'd988, -32'd5842, -32'd1704},
{-32'd5075, -32'd392, 32'd478, 32'd2104},
{-32'd3858, -32'd1777, 32'd4241, -32'd1866},
{32'd2811, 32'd3823, 32'd1805, 32'd4350},
{-32'd11493, 32'd6495, 32'd3647, 32'd984},
{32'd13773, -32'd4098, 32'd1734, 32'd7845},
{32'd4366, 32'd13040, -32'd3115, 32'd5030},
{-32'd4169, -32'd8065, -32'd1440, -32'd4465},
{32'd1782, -32'd9410, 32'd6822, -32'd6836},
{-32'd8387, 32'd8030, 32'd4018, -32'd1667},
{-32'd1878, 32'd268, -32'd6427, -32'd12224},
{-32'd5881, 32'd4570, 32'd2675, 32'd612},
{32'd4079, -32'd4215, 32'd780, 32'd1795},
{32'd3901, 32'd552, 32'd2663, -32'd326},
{-32'd2960, -32'd7372, -32'd7924, -32'd13350},
{-32'd5973, 32'd5759, -32'd1643, -32'd5497},
{-32'd8, -32'd7435, 32'd2769, -32'd273},
{32'd5644, -32'd6387, -32'd10171, -32'd2553},
{32'd12954, -32'd521, 32'd2913, -32'd8215},
{32'd12519, 32'd5525, -32'd5181, 32'd10433},
{32'd8307, -32'd2462, -32'd11554, -32'd973},
{-32'd3703, -32'd7862, 32'd5351, -32'd6308},
{32'd2611, -32'd7168, 32'd6990, 32'd606},
{32'd4926, -32'd3243, 32'd1843, -32'd3205},
{32'd1293, -32'd4176, -32'd24, -32'd3269},
{-32'd247, -32'd3127, 32'd5283, -32'd1021},
{-32'd42, 32'd3953, 32'd344, 32'd5946},
{32'd1468, 32'd2299, 32'd1726, 32'd3512},
{-32'd12128, -32'd4049, -32'd4917, 32'd1949},
{-32'd3213, -32'd1142, 32'd3760, -32'd6732},
{-32'd2347, 32'd1473, 32'd14522, 32'd7415},
{-32'd10736, 32'd1506, 32'd2515, 32'd6061},
{32'd6452, -32'd4261, 32'd2792, 32'd2993},
{-32'd8277, -32'd2176, 32'd3985, -32'd1282},
{-32'd1648, -32'd6990, 32'd10082, -32'd1525},
{32'd6200, -32'd22, 32'd1519, -32'd3364},
{-32'd509, -32'd2151, 32'd405, 32'd2372},
{32'd3376, 32'd2434, 32'd812, -32'd294},
{-32'd3716, 32'd456, -32'd7129, -32'd6599},
{-32'd3569, -32'd9760, -32'd5153, -32'd6898},
{-32'd5, -32'd645, 32'd6659, 32'd4439},
{-32'd7059, -32'd7772, 32'd6283, 32'd7336},
{32'd4962, 32'd1521, -32'd3721, 32'd5143},
{-32'd3342, -32'd1322, -32'd6917, 32'd2127},
{-32'd8548, 32'd104, -32'd2571, 32'd595},
{-32'd9987, 32'd5023, 32'd2685, 32'd246},
{32'd9307, -32'd13717, -32'd3654, -32'd9478},
{32'd2308, 32'd1480, -32'd5320, -32'd40},
{-32'd7787, -32'd5109, 32'd11898, 32'd3236},
{32'd944, 32'd5335, 32'd973, 32'd1316},
{-32'd8901, -32'd5080, 32'd9906, -32'd1672},
{-32'd6200, -32'd7913, -32'd9143, 32'd3736},
{32'd9163, -32'd1866, -32'd969, 32'd1507},
{-32'd977, 32'd1154, -32'd6404, -32'd5576},
{-32'd2389, -32'd6960, 32'd5844, 32'd2661},
{-32'd7952, -32'd2413, 32'd5886, 32'd9543},
{-32'd1786, 32'd3175, 32'd17658, 32'd2392},
{32'd1622, -32'd6918, -32'd15980, -32'd7780},
{32'd4507, 32'd3468, -32'd106, 32'd1627},
{-32'd12352, -32'd2362, 32'd1625, -32'd837},
{32'd6599, 32'd4967, 32'd4464, -32'd180},
{32'd11367, -32'd2812, -32'd1777, -32'd1294},
{-32'd10994, 32'd5044, 32'd6591, 32'd5673},
{32'd7749, 32'd8488, 32'd3072, 32'd707},
{-32'd3785, -32'd6239, 32'd7506, 32'd440},
{32'd8047, -32'd2252, 32'd2624, -32'd2300},
{32'd17293, 32'd1932, -32'd3142, 32'd7156},
{-32'd8688, -32'd7811, -32'd11439, -32'd6380},
{32'd1308, 32'd2912, 32'd4204, 32'd5860},
{32'd1918, -32'd5752, -32'd5893, -32'd1232},
{-32'd1438, -32'd1329, -32'd5884, -32'd455},
{-32'd1566, 32'd2035, -32'd595, 32'd5745},
{-32'd6561, -32'd6175, 32'd1602, 32'd1049},
{-32'd16676, 32'd1767, 32'd4605, -32'd1346},
{-32'd6578, -32'd6340, 32'd993, -32'd300},
{-32'd8535, -32'd8226, 32'd2544, -32'd5303},
{32'd2902, -32'd8178, -32'd7810, -32'd3637},
{32'd4935, -32'd8553, -32'd1302, 32'd1229},
{32'd8365, -32'd6145, 32'd3016, 32'd4955},
{32'd6922, 32'd14179, 32'd6138, 32'd4350},
{-32'd6969, -32'd3791, -32'd349, -32'd2354},
{-32'd1992, 32'd1056, 32'd8528, 32'd7344},
{32'd7857, 32'd1733, -32'd6298, -32'd4601},
{-32'd18233, -32'd796, 32'd2640, -32'd2715},
{32'd7270, -32'd1244, -32'd2809, 32'd3895},
{32'd875, 32'd13397, 32'd8381, 32'd6090},
{-32'd5690, -32'd2779, -32'd3574, -32'd1619},
{-32'd7871, 32'd2324, -32'd5059, -32'd3364},
{-32'd85, -32'd1786, -32'd7080, -32'd5990},
{32'd11147, -32'd4265, 32'd5654, 32'd453},
{32'd1513, -32'd4140, -32'd14572, -32'd694},
{-32'd5081, 32'd3831, -32'd4901, -32'd5185},
{32'd9264, 32'd5213, -32'd3821, 32'd5039},
{32'd10207, -32'd367, -32'd2649, 32'd7488},
{32'd488, 32'd2478, -32'd9220, -32'd5223},
{32'd1652, -32'd7425, 32'd1755, 32'd3772},
{-32'd3007, -32'd4095, -32'd180, 32'd2221},
{32'd8767, -32'd8188, -32'd113, 32'd647},
{-32'd4496, 32'd503, 32'd5953, -32'd3071},
{-32'd3225, -32'd2431, 32'd4818, -32'd2733},
{-32'd2303, 32'd4598, 32'd13140, 32'd647},
{-32'd5325, 32'd298, -32'd4692, -32'd4103},
{32'd10357, -32'd4230, 32'd5273, 32'd610},
{-32'd2208, -32'd2882, -32'd2116, -32'd810},
{-32'd584, 32'd3647, -32'd3115, 32'd909},
{32'd666, -32'd8533, -32'd1659, 32'd3318},
{32'd11306, -32'd469, -32'd7386, -32'd6839},
{-32'd3544, -32'd8575, -32'd659, -32'd3582},
{-32'd2289, 32'd2617, 32'd4747, -32'd3150},
{32'd4740, -32'd7475, -32'd8597, 32'd120},
{-32'd4744, -32'd467, 32'd13991, 32'd5404},
{32'd6599, 32'd2454, -32'd14326, -32'd9753},
{-32'd9051, 32'd2476, 32'd9478, 32'd2922},
{32'd1978, 32'd4503, -32'd6832, 32'd3534},
{32'd3078, -32'd196, -32'd7873, -32'd6942},
{32'd2198, -32'd2038, 32'd12173, 32'd7816},
{32'd3759, 32'd6783, 32'd2727, -32'd3895},
{32'd6530, -32'd2275, -32'd18394, -32'd4878},
{32'd11885, 32'd1105, -32'd13766, -32'd8487},
{32'd13927, -32'd6016, -32'd9362, -32'd3942},
{-32'd10589, 32'd1942, 32'd2894, 32'd7047},
{32'd12396, 32'd6472, 32'd5058, 32'd3012},
{-32'd14163, -32'd3741, -32'd171, -32'd7681},
{32'd9744, -32'd1121, -32'd2844, 32'd2483},
{-32'd9731, -32'd6160, 32'd1977, -32'd1448},
{32'd4606, 32'd10084, 32'd5649, -32'd170},
{-32'd3436, 32'd12679, -32'd12755, -32'd2443},
{-32'd1343, -32'd4930, -32'd14807, -32'd9035},
{-32'd5438, -32'd3730, 32'd6101, 32'd4907},
{32'd8335, 32'd1531, 32'd8537, 32'd8644},
{32'd5750, 32'd6966, 32'd1047, -32'd317},
{32'd3097, -32'd7757, 32'd8924, 32'd3126},
{-32'd4699, -32'd14218, -32'd3907, 32'd5999},
{-32'd3352, -32'd1643, 32'd5771, 32'd1619},
{32'd1442, 32'd1712, 32'd6031, -32'd896},
{32'd9257, 32'd826, 32'd1664, 32'd2820},
{-32'd4501, 32'd6360, 32'd1590, -32'd1212},
{32'd4011, -32'd2143, 32'd4786, -32'd4244},
{32'd291, -32'd3904, -32'd2852, -32'd4046},
{32'd10494, 32'd4192, 32'd5177, 32'd4037},
{-32'd1081, 32'd5580, 32'd202, -32'd2173},
{-32'd2409, -32'd6681, -32'd2025, -32'd9833},
{-32'd12734, 32'd4137, -32'd11716, -32'd2445},
{-32'd4428, -32'd1496, -32'd7985, -32'd4723},
{-32'd6199, -32'd5219, -32'd5753, 32'd383},
{-32'd3954, -32'd628, 32'd10597, 32'd3391},
{-32'd7617, -32'd8371, -32'd4481, -32'd3903},
{32'd13289, 32'd10646, -32'd8752, 32'd4384},
{32'd8502, -32'd2611, -32'd4609, 32'd1420},
{-32'd5213, -32'd12032, -32'd2409, -32'd3947},
{32'd490, 32'd3287, -32'd11442, -32'd5124},
{32'd1966, 32'd13968, 32'd1807, 32'd4982},
{32'd2162, -32'd3514, 32'd11015, 32'd8378},
{32'd1623, -32'd5442, -32'd6238, -32'd8026},
{32'd6685, 32'd3633, 32'd6168, -32'd5358},
{-32'd1346, 32'd1087, 32'd12576, 32'd4758},
{-32'd6545, 32'd1285, -32'd1878, -32'd3406},
{32'd2614, -32'd7124, -32'd5196, -32'd4029},
{-32'd2249, -32'd3340, 32'd5992, -32'd1523},
{32'd6805, 32'd6541, -32'd5512, -32'd3861},
{-32'd19512, -32'd2200, -32'd1572, -32'd2194},
{-32'd7151, -32'd6375, 32'd1744, -32'd7750},
{-32'd1914, -32'd1079, 32'd4363, 32'd3330},
{-32'd4419, -32'd4093, 32'd1767, -32'd3264},
{-32'd4502, 32'd2569, -32'd7809, -32'd38},
{-32'd8343, -32'd1292, -32'd7640, -32'd9842},
{32'd5966, 32'd710, -32'd1356, -32'd6430},
{-32'd3382, 32'd90, 32'd6922, 32'd804},
{32'd1142, 32'd2770, -32'd10042, 32'd1137},
{32'd6482, -32'd4861, -32'd7279, -32'd2493},
{-32'd7199, 32'd13, -32'd2244, 32'd4060},
{-32'd11177, -32'd2054, -32'd8225, -32'd501},
{32'd3225, -32'd2237, 32'd6235, 32'd11528},
{32'd742, 32'd4251, -32'd7099, 32'd4360},
{32'd7793, 32'd384, -32'd2695, 32'd5968},
{-32'd4340, -32'd9549, -32'd4796, -32'd3978},
{32'd361, -32'd8164, 32'd3106, 32'd315},
{-32'd829, 32'd1082, 32'd7808, 32'd9261},
{32'd4429, -32'd3266, 32'd4204, 32'd5388},
{-32'd2356, -32'd5309, 32'd438, -32'd8274},
{32'd2113, -32'd5056, -32'd13662, -32'd10475},
{-32'd7052, -32'd4770, -32'd277, -32'd595},
{32'd9965, -32'd5593, -32'd3115, 32'd3707},
{32'd3805, 32'd10105, -32'd1104, 32'd6376},
{-32'd2045, 32'd4874, 32'd11079, 32'd5632},
{-32'd3565, -32'd5773, 32'd4149, -32'd4652},
{-32'd2583, -32'd6036, -32'd626, -32'd6408},
{32'd16233, 32'd3881, -32'd713, 32'd3795},
{32'd1607, 32'd3008, -32'd4780, 32'd8721},
{32'd15428, 32'd2439, -32'd4034, -32'd738},
{-32'd3248, 32'd529, 32'd1326, 32'd7414},
{-32'd1063, -32'd2857, 32'd4174, 32'd209},
{-32'd899, -32'd14540, -32'd2002, -32'd6423},
{32'd2153, 32'd3270, 32'd5211, 32'd6873},
{-32'd2637, -32'd4822, -32'd6543, -32'd8859},
{32'd2040, -32'd10722, -32'd8584, -32'd1502},
{32'd762, 32'd2112, -32'd5028, -32'd6083},
{-32'd9698, 32'd2853, 32'd1062, 32'd5677},
{32'd4280, 32'd8466, 32'd910, 32'd6548},
{32'd9382, -32'd944, -32'd1391, 32'd1225},
{32'd974, -32'd3321, -32'd8033, 32'd716},
{32'd5032, -32'd1602, -32'd2935, -32'd5199},
{32'd4699, 32'd2501, -32'd5733, -32'd5135},
{32'd2208, -32'd7552, -32'd5754, -32'd6417},
{32'd1533, -32'd228, -32'd1454, 32'd1884},
{-32'd2897, 32'd7740, 32'd21424, 32'd9465},
{32'd9811, -32'd428, 32'd3137, 32'd3294}
},
{{32'd4023, 32'd1998, 32'd8829, 32'd5904},
{-32'd386, -32'd5652, 32'd895, -32'd2102},
{-32'd290, 32'd849, -32'd3121, -32'd4925},
{-32'd6899, 32'd12132, -32'd2571, -32'd2070},
{32'd1235, 32'd3437, 32'd7937, -32'd4173},
{32'd2106, 32'd12048, 32'd2776, -32'd3055},
{-32'd8944, 32'd3793, 32'd7985, -32'd2365},
{32'd4269, -32'd10275, -32'd2324, -32'd10662},
{32'd3504, 32'd2636, -32'd2077, 32'd8083},
{32'd9138, -32'd3603, -32'd5444, 32'd3811},
{-32'd7398, -32'd1366, -32'd898, -32'd5085},
{-32'd5919, -32'd1563, 32'd3085, -32'd1594},
{32'd3076, -32'd3365, -32'd1506, 32'd711},
{32'd3498, 32'd1602, -32'd221, 32'd2288},
{-32'd2551, 32'd1475, 32'd170, -32'd1033},
{-32'd6162, -32'd7447, -32'd7964, -32'd312},
{-32'd11073, 32'd4308, 32'd12454, 32'd4328},
{-32'd341, -32'd283, -32'd13224, -32'd5913},
{32'd812, -32'd11256, -32'd896, -32'd6559},
{-32'd1932, -32'd3696, -32'd8501, 32'd3058},
{-32'd2750, 32'd9048, 32'd4300, 32'd178},
{-32'd7792, 32'd3307, -32'd3134, -32'd404},
{-32'd2772, -32'd11058, 32'd15475, -32'd1640},
{32'd11608, -32'd422, -32'd7314, -32'd4230},
{-32'd1293, 32'd2215, 32'd484, -32'd13414},
{-32'd6428, 32'd6202, 32'd1342, 32'd1150},
{32'd1105, 32'd5389, 32'd9574, -32'd6215},
{32'd2778, 32'd15740, 32'd6766, -32'd255},
{32'd15287, -32'd4852, 32'd2587, -32'd4130},
{-32'd4987, 32'd1229, -32'd6949, 32'd4547},
{-32'd5744, -32'd1465, 32'd8444, 32'd1779},
{-32'd9792, 32'd2151, 32'd12775, 32'd3093},
{32'd8384, -32'd6467, 32'd2030, 32'd3943},
{32'd7506, 32'd1167, -32'd7641, -32'd4630},
{32'd2125, 32'd1855, -32'd9321, -32'd3854},
{32'd1743, -32'd2641, -32'd2271, 32'd5634},
{32'd4448, 32'd3895, -32'd9977, 32'd7062},
{32'd1018, 32'd8324, 32'd6573, -32'd487},
{32'd5515, 32'd1733, 32'd5939, -32'd2472},
{32'd2379, -32'd312, -32'd20071, -32'd2022},
{-32'd57, 32'd1182, 32'd2156, -32'd4181},
{32'd1691, -32'd8505, -32'd13295, -32'd4104},
{-32'd7414, -32'd2512, 32'd1127, 32'd6236},
{32'd2369, 32'd4781, 32'd3124, -32'd5313},
{32'd3356, -32'd2518, -32'd10429, -32'd2921},
{32'd5730, 32'd5839, 32'd4709, 32'd2800},
{-32'd2268, -32'd9233, -32'd3704, 32'd3160},
{32'd1948, -32'd7436, -32'd2925, 32'd2004},
{-32'd7020, -32'd601, -32'd3741, -32'd1388},
{-32'd13091, 32'd11104, 32'd16247, -32'd5859},
{32'd2335, 32'd6284, 32'd6949, 32'd4106},
{-32'd6096, -32'd11364, -32'd8538, -32'd7541},
{32'd879, 32'd10573, 32'd8937, 32'd1884},
{32'd7259, -32'd6287, -32'd3503, 32'd3399},
{32'd6167, -32'd8076, -32'd10517, -32'd3600},
{32'd10323, 32'd442, 32'd5557, 32'd9695},
{32'd5611, 32'd4453, -32'd11652, 32'd8029},
{32'd5930, 32'd771, 32'd5997, 32'd6713},
{-32'd1353, -32'd1057, -32'd5925, -32'd10192},
{-32'd7917, 32'd4260, 32'd5235, 32'd279},
{32'd8106, 32'd18619, 32'd7857, 32'd7774},
{32'd4828, 32'd2043, -32'd5787, -32'd9263},
{-32'd4277, 32'd3074, 32'd2636, -32'd5713},
{-32'd3259, 32'd833, 32'd3039, -32'd580},
{-32'd2358, -32'd5344, 32'd2339, -32'd3995},
{32'd72, 32'd7899, -32'd4213, 32'd4945},
{32'd12375, -32'd3989, 32'd11403, -32'd1581},
{32'd3579, -32'd1759, 32'd909, 32'd6408},
{-32'd12928, -32'd4817, 32'd2486, -32'd2755},
{32'd3394, 32'd9433, -32'd14573, -32'd686},
{-32'd6614, 32'd9481, 32'd8091, -32'd3584},
{-32'd548, 32'd6835, -32'd1171, -32'd3491},
{-32'd1772, -32'd10506, 32'd2518, -32'd1562},
{-32'd771, 32'd1441, 32'd7591, 32'd5076},
{32'd1401, 32'd7379, 32'd2823, 32'd9684},
{32'd19653, -32'd8396, -32'd10569, -32'd7350},
{32'd104, -32'd2709, -32'd9458, -32'd9688},
{-32'd2328, -32'd11632, 32'd10574, 32'd1880},
{32'd15070, 32'd3369, -32'd2407, 32'd263},
{-32'd3423, 32'd1046, -32'd11096, -32'd8762},
{32'd12562, 32'd4124, 32'd4807, -32'd1778},
{-32'd6161, -32'd24037, 32'd4619, 32'd2046},
{32'd1777, -32'd7086, -32'd1206, 32'd3633},
{32'd1084, -32'd14012, 32'd5625, -32'd4950},
{32'd1366, -32'd718, -32'd452, -32'd18610},
{-32'd1333, -32'd3470, 32'd6773, -32'd733},
{32'd11792, 32'd12925, -32'd6370, -32'd7519},
{-32'd1286, -32'd2313, -32'd2877, -32'd4543},
{32'd15773, -32'd1546, -32'd9196, -32'd7657},
{-32'd4359, 32'd2219, 32'd3811, -32'd4355},
{32'd2216, -32'd5736, -32'd5875, 32'd2216},
{-32'd9360, 32'd8446, 32'd10639, -32'd8504},
{32'd5205, -32'd13313, -32'd4147, 32'd604},
{-32'd2871, -32'd9487, -32'd6015, -32'd311},
{-32'd4033, 32'd6652, -32'd7991, 32'd457},
{32'd8166, -32'd10349, 32'd3560, -32'd2484},
{32'd247, -32'd6231, -32'd7951, 32'd5955},
{32'd2416, 32'd2635, -32'd23088, 32'd1407},
{32'd5364, 32'd7421, -32'd3045, 32'd670},
{32'd90, -32'd1312, -32'd2803, -32'd4589},
{-32'd3057, -32'd7219, -32'd4132, -32'd1655},
{-32'd4286, -32'd14228, -32'd11114, -32'd814},
{32'd3182, -32'd13448, -32'd13396, 32'd879},
{32'd18625, 32'd6606, 32'd17283, -32'd17647},
{32'd10738, -32'd4536, 32'd2376, -32'd1635},
{-32'd12931, -32'd1009, 32'd3816, 32'd5220},
{-32'd1693, -32'd1689, -32'd7693, 32'd4452},
{32'd2595, -32'd2776, 32'd6448, -32'd8786},
{-32'd361, 32'd17675, 32'd6332, -32'd1106},
{32'd6700, 32'd6916, -32'd361, -32'd1806},
{-32'd510, -32'd3528, -32'd6511, 32'd1907},
{32'd12683, -32'd7333, 32'd2385, -32'd9555},
{-32'd7410, 32'd1276, 32'd1817, 32'd3990},
{32'd6235, 32'd10397, -32'd2048, -32'd208},
{-32'd1990, -32'd3923, -32'd5020, -32'd5493},
{-32'd3085, 32'd4127, 32'd11225, 32'd4353},
{-32'd863, 32'd3406, 32'd2845, -32'd11182},
{32'd1887, 32'd10914, -32'd764, 32'd3658},
{-32'd10870, 32'd12172, 32'd6673, 32'd11010},
{-32'd6667, 32'd8488, 32'd7672, 32'd1961},
{32'd2100, 32'd14671, 32'd7747, -32'd2400},
{-32'd5475, 32'd6042, -32'd4732, 32'd4103},
{32'd5435, -32'd5703, 32'd9369, -32'd246},
{32'd555, 32'd14594, 32'd5309, 32'd11358},
{-32'd10058, -32'd2363, 32'd6276, -32'd10923},
{32'd1521, 32'd21476, -32'd5599, 32'd7860},
{32'd3833, 32'd298, -32'd2140, -32'd9041},
{-32'd7169, -32'd9335, -32'd7214, 32'd13545},
{-32'd4520, -32'd10588, 32'd7757, 32'd1165},
{-32'd5735, -32'd8554, -32'd5601, -32'd7015},
{-32'd4612, 32'd6345, 32'd19931, -32'd4038},
{32'd4830, -32'd2799, -32'd36, -32'd813},
{-32'd2737, -32'd8871, -32'd285, -32'd1965},
{32'd11547, -32'd5231, -32'd321, -32'd2668},
{32'd7528, -32'd719, 32'd5985, 32'd3095},
{-32'd9150, -32'd8468, -32'd2951, 32'd14554},
{32'd13028, -32'd9702, -32'd11103, 32'd3941},
{-32'd659, -32'd9094, -32'd8494, -32'd1917},
{32'd5814, 32'd2009, -32'd1740, 32'd7411},
{-32'd10172, -32'd4910, -32'd8027, -32'd5616},
{-32'd2990, 32'd8588, 32'd8526, 32'd6027},
{-32'd9846, 32'd8798, -32'd9261, -32'd2617},
{-32'd7701, -32'd754, 32'd15314, -32'd1867},
{-32'd4573, -32'd6648, 32'd10352, -32'd854},
{32'd7003, 32'd1987, -32'd2707, -32'd3681},
{-32'd7220, 32'd3580, 32'd507, 32'd9623},
{-32'd9174, -32'd10446, -32'd5623, -32'd7127},
{32'd9412, 32'd1513, 32'd589, -32'd538},
{-32'd3339, 32'd10448, -32'd7742, 32'd1636},
{-32'd2205, 32'd3991, 32'd3966, -32'd6605},
{-32'd2185, -32'd9878, -32'd5497, -32'd4283},
{32'd3911, -32'd4576, 32'd5375, 32'd18072},
{32'd965, 32'd10601, 32'd9396, 32'd9560},
{32'd10169, 32'd3349, -32'd20738, -32'd9775},
{32'd6095, 32'd6022, -32'd8884, 32'd1877},
{-32'd10648, -32'd1593, -32'd3008, 32'd11201},
{-32'd1021, -32'd7496, -32'd4314, -32'd874},
{32'd13962, -32'd6479, -32'd9644, 32'd940},
{-32'd2851, -32'd13256, 32'd5504, -32'd2630},
{32'd5794, -32'd3945, -32'd12233, 32'd7136},
{32'd3339, 32'd9953, 32'd20454, 32'd380},
{32'd3755, -32'd351, -32'd3230, 32'd276},
{-32'd8005, 32'd16132, 32'd10493, -32'd1288},
{-32'd2409, -32'd5681, 32'd3193, 32'd4885},
{-32'd5264, -32'd5358, -32'd7130, 32'd326},
{32'd2399, -32'd6468, 32'd9305, 32'd2796},
{32'd1093, 32'd6837, -32'd1611, 32'd7043},
{-32'd462, 32'd646, 32'd2600, 32'd4402},
{-32'd2843, -32'd14209, -32'd3170, -32'd6194},
{-32'd4802, 32'd1636, 32'd13388, -32'd7350},
{32'd9379, 32'd3391, -32'd8373, -32'd2607},
{32'd3760, 32'd987, -32'd12905, 32'd3794},
{-32'd1135, -32'd7863, -32'd6271, 32'd4729},
{32'd5712, -32'd14171, 32'd1015, -32'd5536},
{32'd3079, 32'd3334, 32'd1817, 32'd5812},
{32'd1841, -32'd3993, -32'd4906, -32'd8656},
{32'd12867, -32'd5545, -32'd1603, -32'd3948},
{32'd8891, -32'd11799, 32'd1179, 32'd7694},
{-32'd8026, 32'd3074, 32'd6455, -32'd608},
{-32'd10507, 32'd2859, 32'd9861, 32'd1257},
{-32'd6111, -32'd11028, 32'd4947, -32'd1200},
{32'd6266, -32'd15750, 32'd9466, -32'd3788},
{-32'd9856, -32'd8965, 32'd15786, 32'd2189},
{-32'd1532, -32'd6069, -32'd6545, -32'd5455},
{-32'd3475, -32'd2709, -32'd10119, -32'd12814},
{-32'd7601, 32'd6792, 32'd15856, 32'd10732},
{32'd2505, -32'd3805, 32'd4500, 32'd3375},
{32'd72, 32'd1933, 32'd9147, -32'd2216},
{32'd17375, -32'd4244, 32'd1385, 32'd6479},
{-32'd13636, 32'd66, -32'd6401, -32'd1927},
{32'd15054, -32'd2446, -32'd8527, 32'd5482},
{32'd638, 32'd8273, 32'd10323, 32'd3911},
{32'd5370, 32'd912, -32'd946, 32'd940},
{32'd10330, -32'd1817, -32'd6394, -32'd677},
{-32'd10526, -32'd14184, 32'd957, -32'd2206},
{-32'd12797, -32'd2754, 32'd4064, -32'd1735},
{-32'd9942, 32'd2125, 32'd14188, -32'd7067},
{-32'd3509, 32'd4319, 32'd14473, 32'd2451},
{-32'd1751, -32'd11815, -32'd13921, 32'd9501},
{-32'd7115, -32'd8882, -32'd8208, 32'd1859},
{-32'd11862, 32'd2677, 32'd5168, -32'd2020},
{-32'd2171, 32'd5370, -32'd3960, 32'd391},
{-32'd3043, 32'd8090, 32'd3430, -32'd1517},
{32'd1982, 32'd12840, 32'd15661, 32'd13558},
{-32'd1495, -32'd15487, 32'd6683, 32'd2024},
{-32'd252, -32'd2494, -32'd2512, 32'd5650},
{-32'd936, -32'd12843, 32'd12528, 32'd4278},
{-32'd780, 32'd2659, 32'd4371, -32'd1693},
{-32'd3004, 32'd3141, 32'd9040, 32'd2108},
{32'd3519, 32'd1584, -32'd17895, -32'd3250},
{-32'd5050, -32'd4886, -32'd2611, -32'd9275},
{-32'd5903, 32'd3773, 32'd5903, -32'd11047},
{-32'd2525, -32'd2178, 32'd4439, 32'd2966},
{-32'd9205, -32'd5835, 32'd5295, 32'd9553},
{-32'd4441, 32'd2283, 32'd1274, 32'd2554},
{32'd39, 32'd3571, -32'd3994, -32'd9106},
{32'd2804, 32'd13172, -32'd3728, 32'd8070},
{32'd7745, 32'd5618, 32'd7683, -32'd1862},
{32'd4517, -32'd1070, -32'd7677, 32'd5354},
{-32'd8214, 32'd2089, -32'd8167, 32'd6447},
{-32'd2558, 32'd3229, 32'd13392, 32'd655},
{32'd7280, 32'd6443, -32'd4408, -32'd3333},
{32'd5000, 32'd12518, 32'd3473, 32'd1836},
{-32'd2387, 32'd7302, 32'd40, -32'd2258},
{32'd10708, -32'd4545, -32'd916, -32'd4599},
{-32'd4769, 32'd10279, -32'd4589, -32'd912},
{32'd15185, -32'd3765, 32'd1989, 32'd11591},
{32'd1187, 32'd1807, 32'd3743, -32'd3704},
{-32'd1248, -32'd158, 32'd2957, -32'd306},
{-32'd3357, 32'd8653, -32'd1936, 32'd7782},
{-32'd7163, -32'd4389, 32'd1652, -32'd7035},
{32'd11797, 32'd19256, 32'd4194, -32'd5186},
{-32'd10426, 32'd4104, 32'd4349, 32'd9928},
{-32'd2451, -32'd7636, -32'd71, -32'd6000},
{32'd15871, -32'd9507, -32'd6559, -32'd281},
{32'd6407, 32'd6976, -32'd18, 32'd7786},
{32'd10517, 32'd3136, 32'd417, -32'd9775},
{-32'd191, -32'd5653, 32'd9235, -32'd6243},
{32'd556, 32'd9001, 32'd1913, 32'd1172},
{32'd8183, 32'd2920, -32'd9698, -32'd5538},
{-32'd2603, 32'd10815, -32'd4565, 32'd1624},
{-32'd11340, 32'd3203, -32'd145, -32'd4382},
{32'd763, 32'd9363, 32'd9892, -32'd1676},
{-32'd2474, 32'd520, 32'd8238, 32'd6454},
{32'd3988, -32'd7731, -32'd8735, -32'd6247},
{-32'd2843, -32'd12384, 32'd3342, -32'd820},
{32'd6417, -32'd12169, -32'd9346, -32'd2148},
{32'd8993, -32'd4278, -32'd14262, 32'd4187},
{-32'd6228, -32'd399, -32'd11393, -32'd3205},
{32'd5122, 32'd8323, 32'd1162, -32'd4273},
{32'd8976, 32'd6122, 32'd40, -32'd688},
{-32'd1012, -32'd6709, -32'd9880, -32'd6687},
{-32'd5268, 32'd7085, -32'd2188, 32'd14608},
{-32'd1937, 32'd1417, 32'd8755, 32'd2879},
{-32'd6771, 32'd1545, 32'd15381, 32'd5982},
{32'd5891, -32'd1513, -32'd2271, 32'd6326},
{32'd8450, -32'd17028, 32'd993, -32'd2233},
{32'd2805, 32'd5110, 32'd6308, -32'd11740},
{32'd1252, -32'd9938, -32'd5055, -32'd3761},
{32'd2025, 32'd7413, 32'd1569, 32'd6691},
{-32'd11976, 32'd108, -32'd904, 32'd8079},
{32'd5514, -32'd6829, -32'd7856, -32'd2501},
{32'd8501, -32'd11308, -32'd12339, -32'd6486},
{-32'd3065, -32'd5453, -32'd8059, 32'd2265},
{32'd1131, 32'd3197, 32'd10112, 32'd4995},
{-32'd16026, 32'd4431, -32'd4637, 32'd2725},
{32'd7928, -32'd2044, -32'd8092, -32'd372},
{-32'd7999, 32'd8068, 32'd894, -32'd1487},
{-32'd4800, -32'd9289, -32'd13232, -32'd2359},
{-32'd6849, -32'd4021, 32'd8246, 32'd5098},
{-32'd7311, 32'd2333, 32'd13548, 32'd2499},
{-32'd5008, 32'd3269, 32'd15416, 32'd2835},
{-32'd1972, 32'd4891, 32'd13625, 32'd4762},
{-32'd9602, -32'd6063, -32'd6602, -32'd2582},
{-32'd3724, 32'd6804, 32'd2947, 32'd40},
{32'd2325, -32'd699, -32'd1155, 32'd838},
{32'd2610, 32'd924, -32'd6346, 32'd2712},
{-32'd1010, -32'd1839, 32'd4183, -32'd1190},
{32'd2662, 32'd8080, 32'd2097, 32'd3957},
{32'd2383, -32'd8090, 32'd3863, -32'd2493},
{32'd143, 32'd7740, -32'd3312, 32'd10415},
{-32'd3229, 32'd2690, -32'd2244, 32'd5358},
{-32'd4806, 32'd6047, 32'd6746, 32'd2668},
{32'd363, -32'd4628, 32'd2262, -32'd1436},
{-32'd3265, 32'd1327, -32'd1642, -32'd748},
{-32'd4208, -32'd13061, -32'd2917, 32'd190},
{-32'd3640, 32'd18526, 32'd13598, 32'd5770},
{-32'd12773, 32'd10794, 32'd9364, -32'd1101},
{32'd9928, -32'd7580, -32'd4720, -32'd1424},
{32'd8864, -32'd10499, -32'd6140, 32'd1381},
{-32'd4147, 32'd1176, -32'd3620, 32'd4344},
{32'd10399, -32'd4799, 32'd2572, -32'd1255},
{32'd188, -32'd2353, 32'd1235, 32'd8050},
{32'd2266, -32'd2333, -32'd9716, -32'd10331},
{-32'd6006, 32'd8176, -32'd2247, -32'd862},
{-32'd1175, 32'd1693, -32'd16078, -32'd1548},
{-32'd805, 32'd10499, -32'd14288, -32'd1351},
{32'd9838, 32'd5831, -32'd6564, -32'd9286},
{-32'd11367, -32'd1212, 32'd10473, 32'd3996},
{-32'd1571, -32'd7686, 32'd14451, -32'd4263}
},
{{32'd4367, 32'd7742, 32'd11329, 32'd487},
{-32'd1944, -32'd8775, 32'd1563, -32'd8821},
{-32'd8928, 32'd519, -32'd1204, 32'd6682},
{-32'd9637, -32'd1906, -32'd5852, 32'd2924},
{32'd2349, 32'd6223, -32'd793, 32'd7167},
{-32'd477, 32'd5527, -32'd450, -32'd7799},
{32'd10519, 32'd2655, 32'd7589, 32'd13235},
{-32'd405, -32'd12199, -32'd4539, 32'd7849},
{-32'd3315, 32'd914, 32'd690, 32'd1368},
{32'd5797, 32'd3080, 32'd3358, -32'd2856},
{32'd6059, 32'd3373, 32'd4011, -32'd9813},
{-32'd243, -32'd18326, 32'd17606, -32'd8677},
{32'd4340, -32'd4311, -32'd16665, -32'd6811},
{32'd3574, -32'd13822, -32'd5100, 32'd8606},
{-32'd15062, -32'd6432, -32'd196, -32'd8445},
{-32'd15602, -32'd752, -32'd8499, -32'd326},
{-32'd10719, 32'd3097, 32'd10013, 32'd10738},
{-32'd15849, 32'd13211, -32'd4417, -32'd3360},
{32'd268, -32'd8721, 32'd6102, 32'd1859},
{-32'd1761, -32'd415, 32'd7569, 32'd7722},
{32'd74, -32'd9299, 32'd3990, -32'd5120},
{-32'd3009, -32'd3857, 32'd199, -32'd746},
{-32'd6348, -32'd4763, 32'd2246, -32'd965},
{-32'd10878, 32'd6725, 32'd1330, 32'd1878},
{32'd11334, 32'd7689, 32'd1629, -32'd7814},
{-32'd3384, 32'd4720, 32'd11934, 32'd3233},
{-32'd7613, -32'd86, -32'd16424, 32'd3436},
{32'd4696, 32'd3001, -32'd704, -32'd936},
{32'd999, 32'd8372, 32'd1293, 32'd7056},
{32'd4495, 32'd1761, -32'd1516, 32'd7483},
{-32'd10084, 32'd1623, 32'd1074, 32'd4466},
{-32'd7109, 32'd4007, -32'd6043, 32'd6490},
{32'd5982, 32'd7356, 32'd180, 32'd1519},
{-32'd1362, -32'd3748, -32'd3385, -32'd7111},
{32'd1802, 32'd1726, 32'd5314, -32'd679},
{32'd891, -32'd4396, -32'd6824, -32'd5018},
{32'd7948, 32'd6439, 32'd9381, 32'd17153},
{32'd6730, -32'd5883, 32'd15064, -32'd12875},
{-32'd2605, 32'd8581, 32'd11167, -32'd1154},
{-32'd2552, 32'd7240, 32'd9176, -32'd13317},
{-32'd17980, -32'd3935, -32'd3357, -32'd13677},
{-32'd5639, -32'd6258, -32'd2790, -32'd3278},
{32'd7679, -32'd5211, 32'd1815, -32'd4624},
{32'd3878, -32'd9419, 32'd2635, -32'd11321},
{-32'd4353, -32'd945, -32'd10066, -32'd8119},
{32'd2105, -32'd3089, 32'd1899, -32'd6094},
{32'd3501, -32'd7497, -32'd19157, -32'd868},
{-32'd15691, -32'd3611, -32'd12629, 32'd6842},
{32'd7495, 32'd9111, 32'd5417, 32'd7672},
{-32'd4929, 32'd6476, 32'd6047, -32'd3072},
{-32'd8718, 32'd5565, -32'd11828, 32'd2519},
{32'd5213, 32'd45, 32'd4287, -32'd14236},
{32'd8796, -32'd13470, -32'd2526, 32'd9887},
{-32'd6989, -32'd2542, -32'd2822, -32'd11358},
{32'd7569, 32'd968, -32'd10415, -32'd1374},
{-32'd244, -32'd3707, 32'd6135, -32'd3812},
{32'd7793, -32'd5622, 32'd17081, 32'd11335},
{-32'd4335, 32'd7754, 32'd247, 32'd4141},
{-32'd3183, -32'd11695, 32'd2490, -32'd3271},
{32'd4548, -32'd7210, 32'd10375, 32'd240},
{-32'd3860, -32'd5403, 32'd1248, 32'd4018},
{32'd3026, 32'd1715, -32'd10588, 32'd4715},
{-32'd14740, 32'd2050, -32'd5016, 32'd9161},
{-32'd8105, -32'd10769, -32'd3971, 32'd7399},
{32'd6404, -32'd5312, 32'd5166, -32'd8041},
{32'd22764, 32'd1952, 32'd3679, -32'd1253},
{32'd2468, -32'd9146, 32'd13558, 32'd2570},
{-32'd4714, 32'd4645, 32'd2264, 32'd913},
{-32'd12226, -32'd5928, -32'd6348, -32'd6147},
{-32'd1725, -32'd4901, -32'd369, 32'd8893},
{-32'd470, 32'd5481, -32'd2380, -32'd946},
{32'd7746, 32'd4386, 32'd2631, -32'd6575},
{-32'd10649, 32'd6914, -32'd6618, -32'd3466},
{-32'd6890, -32'd3411, -32'd621, 32'd472},
{32'd10460, 32'd7415, 32'd14064, 32'd18413},
{-32'd7109, 32'd9105, 32'd242, 32'd2432},
{-32'd13849, -32'd6289, 32'd1921, -32'd5731},
{-32'd4707, -32'd7487, -32'd1474, 32'd9049},
{32'd10610, -32'd2967, -32'd3361, 32'd5514},
{-32'd18284, -32'd6556, 32'd7916, -32'd2357},
{32'd6147, 32'd2263, 32'd4468, 32'd5267},
{-32'd13235, -32'd15461, -32'd1337, -32'd8486},
{-32'd7259, 32'd244, -32'd6435, 32'd3775},
{32'd7989, 32'd3465, 32'd8399, -32'd5006},
{-32'd54, 32'd9650, -32'd9154, -32'd9100},
{32'd7835, 32'd1693, 32'd6952, -32'd6236},
{32'd2356, 32'd5024, 32'd719, -32'd518},
{-32'd8714, 32'd3212, 32'd5934, -32'd8978},
{-32'd10653, 32'd7, 32'd6413, -32'd4615},
{-32'd10216, -32'd7554, -32'd2586, 32'd10811},
{32'd7228, 32'd1441, -32'd1392, -32'd5098},
{32'd4915, 32'd44, 32'd1793, 32'd1881},
{32'd7343, 32'd4773, -32'd5310, -32'd9829},
{32'd17159, -32'd1609, 32'd4871, 32'd1793},
{32'd417, 32'd14622, -32'd1346, 32'd990},
{32'd985, 32'd10181, -32'd10585, 32'd5666},
{32'd573, 32'd695, 32'd4791, -32'd1096},
{32'd5736, 32'd11526, -32'd8289, 32'd483},
{-32'd939, 32'd3434, -32'd6147, 32'd2882},
{32'd1367, 32'd7599, 32'd4950, -32'd2278},
{-32'd4028, -32'd4656, 32'd9067, -32'd2159},
{-32'd11025, -32'd3859, 32'd4757, -32'd6284},
{-32'd4218, -32'd2904, 32'd4154, -32'd2092},
{-32'd3353, -32'd12857, 32'd3497, -32'd2423},
{-32'd2681, -32'd5173, 32'd1657, -32'd13186},
{32'd4370, 32'd2984, -32'd7383, 32'd13854},
{-32'd3475, 32'd2767, -32'd9419, 32'd147},
{32'd1131, -32'd922, -32'd1728, -32'd5984},
{-32'd6194, -32'd6575, -32'd5430, -32'd2786},
{-32'd6669, 32'd356, -32'd2080, -32'd3032},
{-32'd3235, 32'd7444, -32'd2233, -32'd4492},
{-32'd3241, -32'd6021, 32'd9161, -32'd5878},
{32'd13183, 32'd2020, 32'd1334, 32'd8129},
{32'd1368, -32'd2291, -32'd3144, -32'd7312},
{32'd3364, -32'd305, -32'd7737, -32'd1331},
{-32'd415, -32'd651, -32'd11421, 32'd16079},
{32'd9983, 32'd15385, 32'd9315, 32'd8497},
{32'd9422, 32'd4706, -32'd1034, 32'd5683},
{-32'd2776, 32'd6289, 32'd3841, 32'd246},
{32'd7323, 32'd1872, 32'd5327, -32'd3301},
{-32'd2134, 32'd1624, -32'd4134, -32'd6754},
{32'd6900, -32'd5363, 32'd5205, -32'd4038},
{32'd2855, -32'd6305, 32'd2811, -32'd2386},
{-32'd4898, 32'd2955, 32'd1136, 32'd9921},
{32'd3279, -32'd11861, 32'd251, 32'd10930},
{-32'd3817, 32'd5463, -32'd6100, 32'd20728},
{-32'd1391, 32'd406, -32'd9171, -32'd7409},
{32'd2362, 32'd7334, 32'd9473, 32'd5026},
{-32'd7990, -32'd11651, 32'd7549, 32'd8488},
{-32'd3888, 32'd3314, -32'd345, 32'd1074},
{-32'd2751, 32'd219, -32'd11504, -32'd11471},
{32'd330, 32'd557, 32'd1528, -32'd1545},
{32'd3836, -32'd7718, -32'd6809, 32'd3814},
{32'd9095, 32'd479, 32'd2668, 32'd8093},
{-32'd10981, 32'd5648, -32'd7418, 32'd155},
{32'd1949, 32'd10205, -32'd2188, -32'd1617},
{32'd7109, 32'd1353, -32'd5641, 32'd628},
{-32'd2948, -32'd2361, -32'd13930, -32'd13311},
{-32'd3660, -32'd940, 32'd2532, 32'd5046},
{-32'd12963, -32'd1774, -32'd10023, 32'd1378},
{-32'd7464, -32'd3335, 32'd717, 32'd543},
{-32'd12002, -32'd6356, 32'd5885, 32'd3601},
{32'd3493, 32'd16600, -32'd6159, -32'd1210},
{-32'd5805, 32'd1810, -32'd12169, 32'd11532},
{32'd5694, -32'd3641, 32'd1451, -32'd4287},
{32'd1481, 32'd20096, -32'd1209, 32'd5462},
{-32'd9273, -32'd8488, 32'd4863, -32'd7973},
{-32'd2131, 32'd9530, -32'd5153, -32'd628},
{-32'd7233, 32'd10473, 32'd2099, 32'd5172},
{32'd527, -32'd5733, -32'd10979, -32'd4597},
{-32'd2139, 32'd6608, -32'd8231, 32'd3159},
{32'd4543, -32'd7226, -32'd2916, -32'd449},
{-32'd3067, -32'd8581, -32'd9826, -32'd4877},
{-32'd3858, 32'd8307, -32'd2742, 32'd587},
{-32'd7281, 32'd6577, -32'd7496, 32'd5328},
{32'd4860, 32'd2253, -32'd2533, 32'd11829},
{-32'd5793, -32'd6790, -32'd1539, -32'd3050},
{32'd558, 32'd601, -32'd1575, 32'd1715},
{-32'd8652, -32'd7100, 32'd1936, 32'd5626},
{32'd82, -32'd6122, -32'd13542, 32'd4497},
{32'd832, -32'd7327, -32'd14851, 32'd1247},
{32'd10059, -32'd4689, 32'd3075, 32'd3645},
{-32'd4299, 32'd9049, -32'd19881, -32'd14335},
{32'd6286, 32'd4247, 32'd16092, -32'd2599},
{32'd788, 32'd8457, -32'd4379, -32'd6035},
{-32'd128, -32'd3003, -32'd7393, -32'd11995},
{32'd9507, 32'd14898, -32'd198, 32'd6891},
{-32'd2978, -32'd4182, 32'd1811, -32'd1070},
{32'd4795, -32'd1416, -32'd7459, 32'd2775},
{32'd4355, -32'd9939, 32'd8229, 32'd6007},
{-32'd1248, -32'd8097, 32'd1498, 32'd157},
{32'd12265, 32'd5799, 32'd6991, 32'd20721},
{32'd1658, 32'd408, 32'd6667, 32'd2454},
{32'd3678, 32'd4463, -32'd3340, -32'd4127},
{32'd2217, -32'd5632, -32'd3053, 32'd3159},
{32'd7865, -32'd15184, -32'd5320, -32'd3425},
{-32'd9791, -32'd4821, 32'd3820, 32'd3511},
{32'd302, 32'd6168, 32'd7732, 32'd4913},
{32'd11236, 32'd216, 32'd11072, -32'd7680},
{-32'd6801, 32'd9911, 32'd3401, 32'd3947},
{-32'd6513, 32'd5647, -32'd1171, 32'd2087},
{-32'd18855, -32'd3305, -32'd12299, -32'd5786},
{-32'd732, -32'd3517, -32'd7404, -32'd4959},
{32'd4290, 32'd1981, -32'd9844, 32'd5201},
{32'd3305, 32'd1634, 32'd692, -32'd6578},
{-32'd5689, 32'd2710, -32'd5807, -32'd5253},
{32'd11291, -32'd6589, -32'd10743, 32'd3990},
{-32'd7516, 32'd11913, 32'd5905, 32'd3800},
{32'd4897, 32'd3142, 32'd10221, 32'd5728},
{-32'd5143, 32'd6470, 32'd5382, -32'd7354},
{32'd9464, 32'd1911, -32'd7053, 32'd2452},
{-32'd299, -32'd5550, -32'd14497, -32'd11330},
{-32'd20102, 32'd6571, 32'd8261, 32'd3297},
{32'd3320, 32'd5593, 32'd1366, 32'd2959},
{-32'd11767, 32'd5690, -32'd1191, 32'd15683},
{-32'd3334, -32'd5403, -32'd8368, -32'd2997},
{-32'd11644, 32'd1443, 32'd1424, -32'd3434},
{-32'd1150, 32'd5361, -32'd4019, -32'd6752},
{-32'd9074, 32'd12917, -32'd5267, 32'd3748},
{32'd7781, 32'd683, -32'd13200, 32'd1548},
{-32'd1698, -32'd3952, -32'd8712, 32'd2352},
{32'd7555, 32'd7218, 32'd6653, -32'd15060},
{-32'd8662, 32'd2363, -32'd4276, -32'd3380},
{32'd7004, -32'd9636, 32'd5974, 32'd16931},
{32'd1782, -32'd4819, 32'd2132, -32'd8520},
{32'd4475, -32'd5673, 32'd10991, 32'd1056},
{32'd2486, 32'd2966, 32'd3470, 32'd4986},
{-32'd6964, 32'd899, 32'd957, -32'd7313},
{32'd100, -32'd2481, -32'd7526, 32'd18428},
{-32'd4318, 32'd2398, -32'd5343, -32'd6325},
{-32'd3668, -32'd7767, 32'd280, -32'd5804},
{32'd2942, 32'd1941, 32'd921, -32'd3519},
{-32'd2677, 32'd10626, 32'd8800, -32'd2870},
{-32'd9071, 32'd842, 32'd2336, 32'd2309},
{32'd10312, -32'd3839, -32'd5193, -32'd4175},
{-32'd6303, -32'd4333, 32'd6751, 32'd1727},
{-32'd156, 32'd2489, -32'd2192, 32'd20795},
{-32'd6294, 32'd4476, 32'd2504, -32'd1966},
{32'd7680, -32'd2738, 32'd10483, 32'd15382},
{32'd3007, 32'd6384, -32'd3179, 32'd739},
{-32'd3909, 32'd8129, 32'd4007, 32'd2196},
{-32'd6969, 32'd7038, -32'd1773, -32'd6188},
{32'd2029, 32'd3354, -32'd2895, 32'd13863},
{-32'd5058, 32'd4964, -32'd8633, -32'd2124},
{32'd2405, -32'd4164, -32'd5365, -32'd13390},
{32'd4683, -32'd5771, -32'd5390, 32'd3034},
{-32'd12391, -32'd1387, 32'd15222, -32'd543},
{-32'd3309, -32'd5876, 32'd8605, 32'd7912},
{-32'd614, 32'd3089, -32'd3432, 32'd1914},
{32'd10593, -32'd4702, -32'd400, 32'd3987},
{-32'd838, -32'd11618, -32'd6945, 32'd2460},
{-32'd10608, 32'd5416, 32'd7534, -32'd3686},
{-32'd9482, 32'd6353, -32'd2524, 32'd5458},
{32'd2022, 32'd4226, -32'd2921, -32'd13152},
{32'd5066, 32'd2929, -32'd10116, -32'd2658},
{-32'd804, 32'd3343, -32'd10008, 32'd309},
{32'd6087, -32'd10001, -32'd2848, -32'd10666},
{-32'd3879, -32'd438, -32'd12147, -32'd3054},
{-32'd1451, -32'd1193, 32'd13846, -32'd1652},
{-32'd328, 32'd3509, -32'd1683, -32'd3564},
{-32'd61, 32'd5953, 32'd6668, 32'd1809},
{32'd7669, 32'd2253, -32'd7477, 32'd3086},
{-32'd10907, 32'd5824, -32'd12062, 32'd5440},
{32'd2299, 32'd14367, 32'd17347, -32'd2418},
{32'd3770, -32'd1683, 32'd5156, -32'd5485},
{-32'd534, -32'd7237, -32'd186, 32'd15014},
{-32'd3183, 32'd4785, -32'd6134, 32'd3729},
{-32'd12046, -32'd577, -32'd2710, 32'd2355},
{-32'd5020, 32'd5447, -32'd431, 32'd7003},
{-32'd14757, 32'd1739, 32'd2073, -32'd3574},
{-32'd6034, -32'd3779, -32'd676, 32'd3288},
{-32'd6517, -32'd2154, -32'd8109, 32'd2389},
{-32'd2799, 32'd9885, 32'd4304, 32'd6722},
{-32'd589, -32'd1999, -32'd4775, -32'd8171},
{-32'd11150, 32'd4605, -32'd731, 32'd1451},
{-32'd1356, 32'd8278, 32'd1187, 32'd8408},
{-32'd13857, -32'd6574, -32'd8759, -32'd7251},
{32'd18159, 32'd11296, -32'd1842, 32'd1352},
{-32'd3464, 32'd353, 32'd5939, -32'd12657},
{32'd9178, -32'd1280, 32'd10482, -32'd2957},
{32'd4962, 32'd5132, 32'd1528, 32'd11166},
{-32'd5932, -32'd1409, -32'd962, -32'd6889},
{-32'd8083, -32'd7950, 32'd1894, 32'd8087},
{32'd7186, 32'd7348, -32'd3899, 32'd1522},
{-32'd2331, 32'd1774, 32'd8828, -32'd1587},
{-32'd3718, 32'd10968, -32'd373, -32'd196},
{32'd7637, 32'd6490, -32'd7246, 32'd8538},
{32'd3350, 32'd7335, -32'd1057, -32'd172},
{-32'd10084, 32'd4581, -32'd3506, -32'd5778},
{32'd2388, -32'd3119, 32'd2640, 32'd8754},
{32'd3975, 32'd4755, 32'd2147, 32'd5995},
{32'd8618, -32'd5948, 32'd7693, 32'd7484},
{-32'd18159, 32'd7500, -32'd1057, 32'd3999},
{-32'd1244, -32'd7672, 32'd5645, 32'd1688},
{-32'd1037, -32'd7728, -32'd4633, -32'd11808},
{32'd937, -32'd8748, 32'd11055, 32'd5380},
{32'd11456, 32'd1289, 32'd4488, -32'd3876},
{-32'd11102, 32'd4825, -32'd1032, 32'd2091},
{-32'd11143, 32'd1608, 32'd7286, 32'd4672},
{32'd2209, -32'd14853, -32'd3999, -32'd5263},
{32'd5340, 32'd3600, 32'd14928, -32'd1406},
{32'd2003, 32'd6098, 32'd3366, 32'd3794},
{32'd1728, -32'd406, 32'd3336, 32'd14083},
{32'd7583, 32'd5221, -32'd2133, 32'd564},
{-32'd629, -32'd4408, 32'd7071, -32'd10452},
{32'd1671, -32'd15050, -32'd5586, 32'd5746},
{32'd7182, 32'd1767, 32'd12020, 32'd7950},
{-32'd2663, 32'd2972, -32'd7876, -32'd5950},
{32'd19153, -32'd3362, -32'd145, -32'd539},
{-32'd512, -32'd5407, 32'd2048, -32'd15686},
{-32'd20126, -32'd6787, -32'd364, 32'd5026},
{32'd10591, -32'd4973, -32'd6278, -32'd7040},
{-32'd9968, 32'd8751, 32'd10551, 32'd1140},
{-32'd4857, -32'd5815, 32'd977, -32'd7881},
{-32'd4750, 32'd16020, -32'd584, -32'd1185},
{32'd5019, 32'd8087, -32'd3405, -32'd2197},
{-32'd6653, 32'd1308, 32'd715, -32'd1608},
{32'd22322, 32'd5870, -32'd1862, -32'd11914},
{32'd9850, -32'd2542, -32'd803, 32'd2874},
{-32'd7919, -32'd10734, 32'd750, -32'd10125}
},
{{32'd4004, 32'd1911, 32'd4171, 32'd11367},
{-32'd9202, -32'd13971, -32'd6545, 32'd2914},
{32'd2321, -32'd3321, 32'd2287, 32'd1717},
{32'd1315, 32'd2439, 32'd3716, -32'd3946},
{32'd174, -32'd4015, 32'd2324, 32'd4743},
{-32'd8363, 32'd3058, -32'd5115, -32'd9486},
{32'd8221, -32'd2812, 32'd1000, 32'd9660},
{32'd3009, -32'd1552, -32'd5465, -32'd1670},
{-32'd1704, 32'd109, 32'd887, -32'd2770},
{32'd10176, 32'd10600, 32'd5125, 32'd4013},
{-32'd8106, -32'd11283, -32'd4146, -32'd4942},
{-32'd5657, -32'd731, 32'd4364, -32'd7323},
{32'd2778, 32'd852, 32'd4827, -32'd4857},
{-32'd13623, 32'd5090, 32'd7199, -32'd5349},
{-32'd3965, 32'd2298, -32'd693, -32'd6712},
{-32'd2683, -32'd5326, 32'd10460, -32'd4729},
{32'd2264, 32'd6666, 32'd7297, 32'd4819},
{-32'd1251, 32'd11765, 32'd7207, -32'd5878},
{-32'd4043, 32'd3598, 32'd1775, 32'd167},
{32'd4068, 32'd6439, 32'd2947, 32'd9260},
{32'd5723, -32'd2560, 32'd1582, -32'd5730},
{-32'd4395, -32'd7632, 32'd3227, 32'd330},
{-32'd565, -32'd7864, -32'd5832, 32'd7517},
{-32'd10258, 32'd2462, -32'd4395, 32'd7265},
{32'd3510, 32'd5512, 32'd949, 32'd2450},
{-32'd1885, -32'd1153, 32'd6263, -32'd4397},
{32'd4880, -32'd140, -32'd56, 32'd4603},
{-32'd4201, 32'd4397, -32'd1385, 32'd8503},
{32'd3770, -32'd659, 32'd6789, 32'd4088},
{-32'd3901, -32'd3077, -32'd5227, -32'd6396},
{-32'd7971, 32'd2698, -32'd1915, -32'd464},
{-32'd4665, -32'd1984, 32'd3286, -32'd8577},
{32'd1924, 32'd2813, 32'd94, -32'd2276},
{-32'd10480, 32'd773, 32'd7216, -32'd7478},
{32'd5678, 32'd10130, 32'd5212, 32'd11025},
{32'd4387, 32'd2416, -32'd4622, 32'd3327},
{-32'd2914, 32'd120, 32'd4394, 32'd2130},
{-32'd2111, -32'd2844, 32'd6513, 32'd4183},
{-32'd3711, 32'd7656, 32'd2977, -32'd1676},
{-32'd3647, 32'd3094, -32'd87, 32'd2790},
{32'd3768, -32'd3361, -32'd2818, 32'd761},
{32'd8504, 32'd5424, 32'd1041, 32'd5312},
{-32'd3644, 32'd8148, 32'd7102, 32'd12247},
{-32'd11930, -32'd12086, 32'd1217, -32'd11597},
{-32'd7643, -32'd5485, -32'd1656, -32'd3880},
{32'd5750, 32'd169, 32'd125, -32'd9682},
{-32'd5454, -32'd12247, -32'd3637, 32'd8154},
{32'd6061, 32'd1254, -32'd15, 32'd187},
{-32'd1775, -32'd3233, 32'd4089, 32'd3944},
{32'd715, 32'd6889, -32'd4137, 32'd935},
{32'd5008, 32'd2878, -32'd3, 32'd5521},
{32'd2652, 32'd695, 32'd2294, -32'd4088},
{32'd211, -32'd3167, 32'd1582, 32'd49},
{-32'd4250, -32'd505, 32'd785, 32'd10234},
{32'd8049, 32'd9341, 32'd9588, -32'd1842},
{32'd2416, -32'd374, -32'd1041, 32'd4256},
{32'd5573, -32'd8321, -32'd1876, 32'd4406},
{32'd6521, -32'd10292, 32'd7594, 32'd9216},
{-32'd7313, -32'd1132, 32'd5192, -32'd9217},
{-32'd3653, 32'd2193, -32'd1475, 32'd7438},
{-32'd268, -32'd1670, -32'd2552, 32'd394},
{-32'd1157, 32'd3401, 32'd2862, -32'd7688},
{-32'd4670, -32'd1440, -32'd2888, 32'd3635},
{32'd2013, -32'd4338, -32'd2864, -32'd3958},
{-32'd154, -32'd7789, -32'd3214, -32'd1000},
{32'd5340, 32'd8601, 32'd2888, 32'd4330},
{32'd4531, -32'd899, -32'd5842, -32'd2969},
{-32'd14717, -32'd185, -32'd5365, 32'd3073},
{32'd9483, 32'd10887, -32'd9831, -32'd7791},
{32'd3265, -32'd2031, -32'd3433, 32'd6856},
{-32'd2213, 32'd1885, -32'd792, 32'd4876},
{-32'd9369, -32'd7109, 32'd4219, 32'd809},
{-32'd9772, -32'd2938, -32'd1855, 32'd0},
{-32'd3609, -32'd7252, -32'd5925, 32'd9513},
{32'd3783, 32'd11905, 32'd264, 32'd2},
{32'd5319, 32'd8175, -32'd16005, 32'd1545},
{-32'd1040, -32'd4037, 32'd3376, -32'd553},
{-32'd1771, 32'd3186, 32'd2632, -32'd1509},
{32'd3260, 32'd4002, 32'd1409, 32'd3414},
{32'd12645, -32'd8010, 32'd7461, 32'd2881},
{-32'd456, 32'd5940, -32'd3219, -32'd3737},
{32'd9379, -32'd689, 32'd3850, 32'd1330},
{32'd3296, -32'd5015, -32'd4210, 32'd4818},
{-32'd31, -32'd1075, 32'd3293, -32'd157},
{32'd4546, -32'd4257, 32'd122, -32'd2280},
{32'd10108, 32'd5477, 32'd243, -32'd7320},
{32'd6643, 32'd2127, 32'd12073, -32'd539},
{-32'd10399, -32'd3902, -32'd419, 32'd3050},
{32'd8981, -32'd561, 32'd704, -32'd3372},
{-32'd3923, 32'd7876, 32'd7565, -32'd1457},
{32'd2269, 32'd7525, 32'd1740, 32'd4375},
{32'd5190, 32'd2452, -32'd8119, -32'd6055},
{-32'd371, 32'd3483, 32'd7294, 32'd2228},
{32'd39, 32'd10592, 32'd4403, 32'd3591},
{32'd1644, 32'd1912, 32'd10771, 32'd1918},
{-32'd10179, -32'd3738, -32'd2030, -32'd14566},
{32'd10767, 32'd6412, 32'd5782, 32'd4611},
{32'd473, 32'd5569, 32'd684, -32'd5478},
{32'd2011, -32'd8435, -32'd4449, -32'd356},
{32'd5534, 32'd10561, 32'd2963, 32'd5206},
{-32'd2451, -32'd2202, 32'd419, -32'd3844},
{-32'd4413, -32'd3979, -32'd5029, -32'd3620},
{-32'd4923, -32'd8579, 32'd1197, 32'd15307},
{32'd13718, -32'd3977, 32'd3728, -32'd5028},
{-32'd5757, -32'd5964, 32'd4717, 32'd15194},
{32'd1493, 32'd2039, -32'd258, -32'd5301},
{32'd1785, -32'd7622, 32'd3948, -32'd1611},
{-32'd1109, 32'd643, 32'd2437, -32'd306},
{32'd5016, 32'd5499, 32'd6310, 32'd6842},
{-32'd11638, -32'd11089, 32'd7305, 32'd9537},
{32'd3606, 32'd1234, -32'd4851, 32'd5060},
{-32'd528, -32'd3050, 32'd1845, 32'd12053},
{32'd7394, -32'd5418, 32'd4843, 32'd3494},
{32'd2584, 32'd6311, -32'd2674, 32'd5606},
{32'd10324, -32'd3255, 32'd3117, -32'd5930},
{-32'd2625, 32'd8627, -32'd8475, 32'd2290},
{32'd4980, -32'd2861, -32'd575, -32'd1978},
{32'd177, 32'd663, -32'd10400, 32'd3928},
{-32'd1857, -32'd1015, -32'd1602, 32'd5547},
{32'd4574, 32'd810, 32'd713, 32'd1765},
{32'd2980, 32'd8255, -32'd2379, -32'd5880},
{-32'd1932, -32'd930, 32'd8128, -32'd1301},
{-32'd6797, -32'd2313, 32'd344, -32'd2299},
{-32'd1558, 32'd290, -32'd7947, 32'd9603},
{-32'd2373, -32'd332, 32'd1130, 32'd762},
{-32'd4158, 32'd4350, -32'd126, -32'd2702},
{32'd864, -32'd837, 32'd8244, -32'd4334},
{-32'd7386, -32'd5579, -32'd7007, 32'd2488},
{-32'd7864, -32'd7514, -32'd2482, -32'd3718},
{-32'd2710, -32'd2125, 32'd4611, 32'd1488},
{32'd6050, 32'd5573, -32'd1513, 32'd13922},
{-32'd6354, -32'd3243, 32'd3180, -32'd2232},
{-32'd6898, 32'd1303, 32'd1802, -32'd4852},
{-32'd7893, -32'd12944, -32'd1089, 32'd13415},
{-32'd12492, 32'd2638, -32'd2062, -32'd5503},
{-32'd8163, 32'd5352, 32'd4953, -32'd2742},
{32'd4694, 32'd2667, -32'd2013, -32'd6881},
{-32'd2535, -32'd6689, -32'd1072, 32'd5477},
{-32'd7282, 32'd4995, -32'd2558, -32'd1595},
{-32'd1800, -32'd1363, -32'd5255, 32'd1982},
{-32'd4972, 32'd2312, -32'd2252, 32'd6046},
{-32'd6916, -32'd4615, 32'd3291, -32'd3034},
{-32'd818, 32'd4812, -32'd5218, 32'd318},
{-32'd7442, 32'd1098, -32'd2746, -32'd37},
{32'd1976, 32'd13701, 32'd3758, 32'd3592},
{-32'd4424, 32'd7794, -32'd1772, 32'd7284},
{-32'd3171, -32'd278, 32'd6900, 32'd1372},
{-32'd1210, 32'd2130, -32'd8915, -32'd1837},
{32'd7384, -32'd2579, -32'd5889, -32'd1266},
{-32'd3008, -32'd4671, -32'd1720, 32'd3459},
{-32'd6671, -32'd3705, 32'd931, -32'd11148},
{32'd6547, 32'd11058, 32'd3109, 32'd5395},
{-32'd6329, 32'd4483, 32'd899, -32'd6149},
{32'd5040, -32'd24, 32'd4513, -32'd8261},
{-32'd9154, -32'd8005, -32'd6318, -32'd2820},
{-32'd2160, -32'd12365, -32'd1917, -32'd202},
{32'd3868, 32'd712, 32'd6006, 32'd10431},
{32'd6326, -32'd2534, -32'd1588, -32'd5574},
{-32'd2286, 32'd5066, 32'd2734, -32'd7902},
{32'd2352, 32'd4454, 32'd1993, 32'd1961},
{-32'd3228, -32'd5645, -32'd1785, 32'd1592},
{32'd9605, 32'd11451, -32'd950, 32'd1974},
{32'd5069, 32'd4922, 32'd1257, 32'd6837},
{-32'd10185, -32'd6002, 32'd2781, -32'd208},
{32'd7948, -32'd170, 32'd3965, 32'd2701},
{-32'd1203, -32'd22, -32'd10152, 32'd7337},
{32'd11033, 32'd1950, -32'd1750, 32'd4564},
{32'd345, -32'd2112, -32'd6998, -32'd6757},
{-32'd5763, -32'd5796, 32'd1027, 32'd2608},
{-32'd5159, -32'd5289, -32'd561, -32'd15394},
{-32'd2743, -32'd7200, 32'd3129, 32'd3938},
{-32'd12328, -32'd8743, -32'd4549, 32'd7744},
{32'd1521, 32'd1, 32'd2881, 32'd8137},
{-32'd629, -32'd2627, 32'd4847, -32'd15996},
{-32'd1592, 32'd4630, 32'd2219, 32'd6809},
{32'd3094, 32'd4289, 32'd3612, -32'd7989},
{32'd731, 32'd736, -32'd4199, -32'd5228},
{32'd7179, -32'd49, -32'd7675, -32'd431},
{-32'd896, -32'd3940, 32'd261, 32'd13068},
{-32'd11472, -32'd5549, 32'd3172, -32'd10417},
{-32'd8623, -32'd2938, 32'd210, 32'd4030},
{-32'd704, -32'd5294, 32'd10879, -32'd11774},
{32'd727, -32'd11518, -32'd5915, 32'd489},
{-32'd3271, 32'd3857, 32'd9588, -32'd7080},
{-32'd7269, -32'd6691, 32'd7518, 32'd5160},
{32'd5518, 32'd6428, 32'd127, -32'd4917},
{32'd2251, 32'd7857, -32'd4748, 32'd8095},
{-32'd1430, 32'd2677, 32'd1299, -32'd8460},
{32'd4655, -32'd13476, 32'd2975, -32'd856},
{-32'd2975, 32'd1434, 32'd953, -32'd7178},
{-32'd1326, -32'd5325, 32'd2029, 32'd4116},
{-32'd11483, -32'd10671, 32'd2249, -32'd4233},
{32'd4656, -32'd478, 32'd7582, 32'd542},
{-32'd295, 32'd4074, 32'd940, -32'd266},
{-32'd4148, -32'd6481, 32'd927, -32'd876},
{-32'd363, 32'd7825, 32'd3908, 32'd4785},
{-32'd344, -32'd3000, -32'd6813, -32'd10035},
{32'd12771, 32'd6757, -32'd1659, -32'd2923},
{32'd1231, -32'd1097, -32'd5438, 32'd8609},
{32'd7111, 32'd476, 32'd99, -32'd8214},
{-32'd9811, -32'd10150, -32'd3359, -32'd4929},
{32'd1518, -32'd602, -32'd1782, 32'd789},
{-32'd8446, -32'd10719, -32'd1006, 32'd7070},
{-32'd2313, 32'd419, -32'd813, 32'd38},
{-32'd438, 32'd903, -32'd4442, -32'd4520},
{32'd2575, -32'd643, 32'd3112, 32'd2158},
{32'd2633, 32'd1382, -32'd950, 32'd7321},
{32'd3801, -32'd152, -32'd4484, -32'd11556},
{-32'd7887, -32'd7163, -32'd34, 32'd7141},
{32'd4011, 32'd5436, 32'd4479, 32'd5214},
{32'd7630, -32'd3735, -32'd7152, -32'd1586},
{32'd6718, 32'd10664, 32'd1512, -32'd7658},
{32'd4619, 32'd1702, -32'd6427, 32'd6874},
{32'd5834, 32'd4912, -32'd1190, -32'd6355},
{-32'd2763, 32'd3829, 32'd36, -32'd2363},
{-32'd4239, -32'd3196, 32'd6311, -32'd1358},
{-32'd4998, 32'd2313, -32'd9177, 32'd2529},
{-32'd2553, -32'd874, -32'd2914, -32'd5851},
{32'd476, 32'd4717, -32'd1213, 32'd1480},
{32'd2706, -32'd3427, -32'd3510, -32'd829},
{-32'd10608, -32'd4589, -32'd3319, -32'd8121},
{32'd6501, -32'd674, -32'd2128, 32'd6802},
{-32'd1799, -32'd7047, 32'd9371, 32'd5548},
{-32'd2079, -32'd9985, 32'd5749, -32'd3420},
{32'd3297, -32'd3898, 32'd1395, -32'd11838},
{-32'd1768, -32'd4757, 32'd5156, 32'd129},
{32'd1170, 32'd6579, -32'd2576, 32'd2187},
{32'd6255, 32'd1201, 32'd1466, -32'd8430},
{-32'd1000, 32'd8378, 32'd5495, 32'd12353},
{32'd7675, -32'd6268, 32'd666, 32'd5374},
{-32'd5140, -32'd1492, -32'd1668, 32'd282},
{-32'd11106, -32'd68, -32'd4132, -32'd7351},
{-32'd1860, 32'd416, -32'd1302, -32'd1382},
{32'd5209, 32'd3818, -32'd4592, -32'd1488},
{-32'd10888, -32'd6304, -32'd10194, -32'd3963},
{32'd5379, -32'd4536, -32'd1035, -32'd871},
{-32'd5877, -32'd2668, -32'd7169, -32'd7072},
{-32'd8715, -32'd4116, 32'd8957, -32'd2333},
{32'd700, 32'd2282, 32'd2232, -32'd9060},
{-32'd2047, -32'd1031, -32'd554, -32'd429},
{-32'd1036, -32'd9384, 32'd4568, -32'd588},
{32'd5910, 32'd10403, -32'd4203, -32'd525},
{-32'd12117, -32'd7048, -32'd4591, -32'd6799},
{32'd3148, -32'd7655, 32'd841, 32'd2748},
{32'd11505, 32'd15092, 32'd5771, -32'd3524},
{-32'd130, -32'd1321, -32'd7170, -32'd2063},
{-32'd3422, -32'd3005, 32'd6459, -32'd844},
{32'd4570, 32'd7152, -32'd904, -32'd540},
{-32'd6094, -32'd6446, 32'd87, -32'd6385},
{32'd432, 32'd3022, -32'd3778, -32'd5596},
{-32'd2559, 32'd5436, -32'd3094, -32'd8514},
{-32'd1470, 32'd4646, 32'd305, -32'd3374},
{-32'd560, 32'd12167, 32'd5310, -32'd1061},
{-32'd9809, -32'd1310, -32'd1415, -32'd1440},
{-32'd7344, -32'd2323, -32'd1718, -32'd816},
{32'd5517, -32'd4913, 32'd5549, 32'd4600},
{32'd382, 32'd94, -32'd2122, 32'd2856},
{32'd4178, 32'd7931, -32'd3560, -32'd11078},
{-32'd602, -32'd164, -32'd269, 32'd782},
{32'd1096, -32'd936, -32'd2777, 32'd899},
{32'd3386, -32'd2290, 32'd360, 32'd4119},
{32'd707, 32'd3399, -32'd358, -32'd5818},
{-32'd8015, -32'd740, -32'd4160, -32'd1549},
{-32'd6638, -32'd6162, 32'd6247, -32'd6457},
{-32'd6067, -32'd6991, -32'd790, 32'd3103},
{-32'd10287, -32'd4863, -32'd1337, -32'd2042},
{-32'd3466, -32'd3377, 32'd6877, -32'd2428},
{-32'd2096, 32'd2519, 32'd8738, 32'd4369},
{-32'd3023, -32'd5287, -32'd2552, 32'd1757},
{32'd2875, 32'd5651, -32'd2604, 32'd8240},
{-32'd6108, 32'd122, -32'd5246, 32'd290},
{32'd93, -32'd10663, -32'd4505, 32'd4004},
{-32'd2923, -32'd636, 32'd1137, 32'd57},
{32'd2308, -32'd4253, -32'd6008, -32'd3410},
{-32'd5941, 32'd3979, 32'd1432, -32'd6718},
{-32'd10800, -32'd5457, -32'd1008, 32'd897},
{32'd13617, 32'd15007, 32'd9040, 32'd127},
{32'd5596, 32'd4623, -32'd4458, -32'd4647},
{-32'd1053, 32'd355, -32'd1388, -32'd14420},
{-32'd2252, -32'd3560, 32'd4421, 32'd796},
{32'd1695, 32'd6709, 32'd2325, 32'd7559},
{-32'd1415, -32'd13155, 32'd3771, 32'd8012},
{-32'd5904, -32'd7870, -32'd2259, 32'd166},
{-32'd1817, -32'd13396, -32'd12428, 32'd4967},
{32'd2767, 32'd1419, 32'd1630, 32'd2650},
{-32'd7664, -32'd4835, -32'd3100, 32'd8483},
{-32'd325, 32'd9562, -32'd3854, 32'd352},
{-32'd6116, -32'd1271, 32'd4948, -32'd2108},
{32'd1198, 32'd7991, 32'd781, -32'd1272},
{-32'd1596, 32'd2046, 32'd6096, 32'd1840},
{-32'd3946, -32'd5798, 32'd2574, -32'd4824},
{32'd9875, 32'd9043, -32'd866, -32'd2427},
{32'd13632, 32'd6797, 32'd5996, 32'd2097},
{-32'd3455, 32'd1876, 32'd188, -32'd5210},
{-32'd2256, -32'd3027, -32'd11786, -32'd1020},
{-32'd960, 32'd863, 32'd958, -32'd9706},
{32'd2604, 32'd1754, 32'd6653, 32'd3114},
{32'd10287, 32'd2078, 32'd4315, 32'd4005},
{-32'd214, -32'd4331, 32'd1028, 32'd12020},
{-32'd6235, 32'd253, 32'd623, 32'd8676}
},
{{32'd5021, 32'd5887, 32'd84, 32'd7708},
{-32'd281, -32'd13311, -32'd3265, -32'd2078},
{-32'd5450, 32'd4017, -32'd369, 32'd1156},
{32'd2003, -32'd8015, 32'd699, 32'd3611},
{32'd14225, 32'd2401, -32'd2083, 32'd1609},
{32'd8915, 32'd7421, 32'd889, -32'd4599},
{-32'd7046, -32'd272, -32'd4828, 32'd4283},
{32'd470, -32'd10621, 32'd1994, -32'd3466},
{-32'd1746, 32'd3928, 32'd6100, -32'd2383},
{32'd9077, 32'd6914, 32'd9316, 32'd6268},
{-32'd3626, 32'd3061, -32'd6889, -32'd4326},
{32'd4787, 32'd4024, 32'd4139, 32'd590},
{32'd5821, -32'd1985, 32'd2328, 32'd180},
{32'd1627, -32'd11452, 32'd1220, 32'd2753},
{-32'd26700, 32'd716, -32'd4642, -32'd2362},
{-32'd3172, -32'd9212, 32'd923, -32'd664},
{32'd12712, 32'd2236, 32'd7467, 32'd1951},
{32'd3173, -32'd5348, 32'd2829, -32'd8746},
{-32'd1329, -32'd2870, -32'd2279, 32'd14671},
{-32'd9360, 32'd1279, -32'd2053, 32'd8179},
{-32'd9225, -32'd16954, 32'd3916, 32'd2548},
{-32'd11170, -32'd5461, -32'd6811, -32'd6183},
{-32'd4588, -32'd1631, -32'd8726, -32'd882},
{-32'd11165, -32'd4560, -32'd3481, -32'd4686},
{32'd70, 32'd11518, 32'd2741, 32'd11586},
{-32'd6721, -32'd8356, -32'd8283, -32'd3622},
{-32'd11207, -32'd151, 32'd1930, -32'd2235},
{32'd6419, 32'd2220, 32'd3737, 32'd2165},
{32'd9882, 32'd2391, 32'd10249, 32'd3367},
{-32'd4470, 32'd6491, -32'd3734, -32'd3817},
{32'd8403, 32'd6479, -32'd11283, -32'd11244},
{-32'd7157, -32'd1087, -32'd3807, -32'd5369},
{32'd1712, 32'd677, -32'd4853, 32'd3936},
{32'd8700, 32'd8636, -32'd1948, -32'd6353},
{32'd4412, 32'd3070, 32'd9438, 32'd5204},
{-32'd9062, 32'd9277, -32'd6757, -32'd2187},
{32'd5428, -32'd8688, 32'd848, 32'd4849},
{-32'd2273, -32'd10774, -32'd1776, 32'd3333},
{32'd488, 32'd3869, 32'd3649, 32'd3471},
{-32'd11654, -32'd803, 32'd5940, -32'd4112},
{32'd1497, -32'd4705, -32'd4458, 32'd4797},
{32'd5226, 32'd566, 32'd2640, 32'd6114},
{32'd9744, 32'd7621, 32'd6461, 32'd50},
{32'd5515, -32'd7609, -32'd836, 32'd3450},
{-32'd11509, 32'd3190, 32'd7851, -32'd6585},
{32'd3835, -32'd2244, 32'd2785, 32'd4158},
{32'd11119, -32'd3438, -32'd8701, -32'd9729},
{-32'd3444, -32'd8002, -32'd1984, -32'd2045},
{-32'd5207, 32'd4047, 32'd4606, 32'd3814},
{-32'd6046, 32'd4859, 32'd8012, 32'd4298},
{32'd13910, -32'd34, 32'd929, -32'd7978},
{-32'd12555, 32'd7236, 32'd4867, 32'd2531},
{32'd1795, -32'd1230, -32'd1872, -32'd6032},
{-32'd6993, -32'd7333, -32'd6477, 32'd8034},
{-32'd3041, -32'd6023, 32'd12839, 32'd2688},
{-32'd1710, -32'd5133, -32'd8594, -32'd3718},
{-32'd415, -32'd2279, 32'd3437, -32'd5002},
{-32'd3805, -32'd183, -32'd9766, 32'd1323},
{-32'd780, -32'd4319, -32'd78, 32'd864},
{32'd2866, 32'd66, -32'd4246, -32'd8138},
{-32'd7379, -32'd7649, 32'd2234, -32'd4676},
{32'd5761, -32'd7120, 32'd5563, -32'd523},
{32'd3689, -32'd5643, -32'd13041, 32'd2469},
{32'd1622, 32'd482, -32'd8202, -32'd2441},
{32'd7136, 32'd11019, -32'd1410, 32'd4183},
{-32'd672, 32'd4753, 32'd6753, -32'd336},
{-32'd956, 32'd5542, -32'd1724, -32'd9560},
{32'd111, -32'd896, 32'd4236, -32'd8783},
{-32'd7334, 32'd13481, 32'd1141, 32'd2824},
{32'd13318, -32'd4146, -32'd1608, 32'd1533},
{-32'd7611, 32'd5453, 32'd3360, 32'd8798},
{32'd1415, -32'd2476, 32'd1142, 32'd2161},
{-32'd15585, 32'd2637, -32'd6083, -32'd2339},
{32'd1773, -32'd523, 32'd6095, -32'd2735},
{-32'd3672, -32'd1452, -32'd3608, -32'd2918},
{-32'd10768, -32'd3675, -32'd1730, 32'd359},
{32'd3384, -32'd9044, 32'd2554, 32'd1458},
{32'd2678, 32'd5297, -32'd4886, 32'd1166},
{-32'd1878, 32'd3770, 32'd6108, 32'd6938},
{-32'd4881, -32'd16332, 32'd2712, 32'd4085},
{-32'd245, -32'd6277, 32'd10982, -32'd1484},
{32'd8991, 32'd3184, 32'd4314, 32'd3693},
{32'd13073, 32'd1762, -32'd950, 32'd3490},
{32'd2304, 32'd1700, 32'd4467, 32'd745},
{32'd9073, -32'd2740, 32'd4999, -32'd4475},
{-32'd2729, 32'd10679, 32'd1396, 32'd7718},
{-32'd11691, -32'd5706, 32'd9692, 32'd9089},
{32'd2551, -32'd10529, -32'd5649, 32'd999},
{32'd5501, 32'd6877, -32'd1070, 32'd5987},
{-32'd2691, -32'd8203, 32'd3273, 32'd6731},
{-32'd2978, 32'd9364, 32'd577, 32'd2052},
{-32'd11858, -32'd5261, -32'd4172, 32'd5335},
{-32'd3537, -32'd4921, -32'd2193, 32'd1725},
{32'd12369, 32'd8368, 32'd6724, 32'd903},
{-32'd387, -32'd896, -32'd1000, 32'd252},
{-32'd4673, -32'd7123, -32'd3774, 32'd6703},
{32'd12523, 32'd10355, 32'd3173, -32'd840},
{32'd5276, 32'd2299, -32'd1185, -32'd5550},
{32'd8723, 32'd10094, 32'd1485, -32'd3962},
{32'd7909, 32'd2957, 32'd8966, 32'd6068},
{-32'd2042, -32'd2390, 32'd10843, -32'd5384},
{32'd3069, 32'd223, -32'd742, -32'd3909},
{32'd9893, -32'd7097, -32'd881, -32'd5587},
{32'd7879, 32'd5333, 32'd4350, 32'd5930},
{32'd8277, -32'd6307, -32'd1143, 32'd2824},
{-32'd10146, -32'd1758, -32'd9360, 32'd3},
{-32'd824, 32'd226, -32'd9485, -32'd5842},
{-32'd5047, 32'd7680, -32'd2122, -32'd11694},
{32'd3030, 32'd2794, 32'd4871, 32'd10054},
{-32'd5178, -32'd3057, -32'd4104, -32'd7400},
{32'd2886, -32'd6765, 32'd5620, -32'd4971},
{32'd12619, 32'd2918, 32'd5148, 32'd8931},
{32'd1116, 32'd14203, -32'd2751, 32'd6019},
{-32'd1995, -32'd3228, -32'd2234, -32'd104},
{-32'd1707, -32'd10588, -32'd3330, 32'd819},
{-32'd1242, -32'd2786, -32'd4605, 32'd4276},
{32'd2430, 32'd9695, 32'd2081, 32'd1932},
{-32'd10408, 32'd9109, 32'd2855, -32'd1850},
{32'd17010, 32'd3935, -32'd5309, -32'd5221},
{32'd4285, 32'd4151, 32'd1267, 32'd4590},
{-32'd5130, -32'd3157, 32'd1236, 32'd5510},
{-32'd4733, -32'd3441, -32'd772, 32'd6492},
{32'd2865, -32'd2299, 32'd4119, 32'd192},
{-32'd5871, 32'd5132, -32'd5181, -32'd4716},
{32'd11327, 32'd308, 32'd3849, 32'd1716},
{32'd6121, -32'd1936, 32'd5715, 32'd3565},
{-32'd9789, -32'd2503, -32'd2237, -32'd3430},
{-32'd4489, -32'd4020, 32'd1994, -32'd659},
{-32'd253, -32'd9323, -32'd6984, -32'd11408},
{-32'd578, -32'd4087, 32'd7071, -32'd158},
{32'd3636, 32'd2052, -32'd5081, 32'd5504},
{-32'd13941, 32'd7785, -32'd4402, -32'd10090},
{-32'd14451, 32'd4333, 32'd1817, -32'd613},
{32'd601, 32'd12616, 32'd5097, 32'd804},
{32'd6237, 32'd7598, -32'd4902, 32'd3901},
{-32'd4233, 32'd2884, -32'd556, -32'd2723},
{32'd1041, -32'd10165, -32'd8029, 32'd6660},
{-32'd6097, -32'd1269, 32'd3932, 32'd2683},
{-32'd3175, -32'd2562, -32'd781, -32'd2261},
{-32'd8735, -32'd2534, -32'd3297, -32'd4831},
{32'd1760, 32'd7231, -32'd654, 32'd7624},
{-32'd1296, 32'd2714, -32'd4710, 32'd559},
{-32'd11005, -32'd5756, -32'd5049, -32'd6270},
{32'd1177, -32'd3917, 32'd1949, 32'd4202},
{32'd19054, 32'd2564, 32'd6847, 32'd1001},
{32'd5862, -32'd405, 32'd6930, -32'd8222},
{-32'd7569, -32'd5555, 32'd4834, -32'd4608},
{-32'd11020, -32'd5785, -32'd14, 32'd1184},
{-32'd5894, -32'd6738, 32'd6028, -32'd609},
{32'd1491, -32'd16159, -32'd119, -32'd6338},
{32'd4589, -32'd1435, -32'd7446, 32'd3933},
{32'd5015, 32'd2303, -32'd1270, 32'd1704},
{32'd9470, -32'd8662, -32'd6388, 32'd1751},
{32'd1990, -32'd6584, -32'd1115, -32'd4529},
{-32'd1446, 32'd3557, -32'd4402, 32'd1055},
{-32'd7869, -32'd6091, -32'd3405, -32'd1732},
{32'd12509, 32'd9336, 32'd4462, 32'd7871},
{32'd13043, -32'd3013, 32'd4624, 32'd1843},
{32'd6219, 32'd5323, -32'd2960, -32'd6538},
{-32'd3500, 32'd7056, -32'd2186, 32'd693},
{-32'd2371, -32'd2075, -32'd2055, 32'd273},
{32'd15590, -32'd2203, -32'd3287, -32'd4315},
{-32'd934, 32'd9897, -32'd4048, -32'd10283},
{32'd15879, 32'd888, 32'd5738, -32'd2734},
{32'd1028, -32'd395, 32'd7437, -32'd13308},
{-32'd17457, -32'd871, -32'd229, 32'd2236},
{-32'd12542, -32'd9542, 32'd3459, -32'd2462},
{-32'd13510, 32'd3066, -32'd170, -32'd2109},
{-32'd1827, 32'd245, -32'd5226, 32'd4354},
{32'd3928, -32'd6398, -32'd6228, 32'd1596},
{-32'd8473, 32'd4728, 32'd2149, -32'd1974},
{-32'd10655, -32'd1298, -32'd3682, -32'd2317},
{32'd7779, 32'd4092, 32'd5333, 32'd3525},
{-32'd5411, -32'd75, -32'd2810, -32'd1170},
{32'd10916, 32'd440, -32'd9690, -32'd3403},
{32'd2437, -32'd1526, -32'd1526, 32'd4529},
{32'd8091, -32'd8465, 32'd12010, -32'd5649},
{32'd2715, -32'd4129, -32'd1868, -32'd3783},
{-32'd854, -32'd8178, -32'd3314, 32'd3150},
{-32'd8926, -32'd11003, -32'd716, -32'd5526},
{-32'd1995, -32'd8170, -32'd10848, -32'd6982},
{-32'd3311, -32'd1103, -32'd2981, 32'd1134},
{32'd3453, 32'd8507, -32'd1743, -32'd8436},
{32'd2059, 32'd6638, 32'd7801, 32'd4044},
{-32'd5022, -32'd1246, -32'd1281, -32'd2168},
{32'd9331, 32'd2125, -32'd836, 32'd4038},
{-32'd4995, 32'd6309, 32'd7334, -32'd3921},
{-32'd4661, -32'd2051, 32'd3030, -32'd12575},
{-32'd9085, 32'd1465, 32'd2245, -32'd4839},
{-32'd1628, -32'd5476, -32'd4261, 32'd1803},
{32'd2270, 32'd917, -32'd3769, 32'd2045},
{-32'd12082, 32'd6366, -32'd3222, -32'd129},
{-32'd4143, -32'd3475, 32'd5826, 32'd936},
{-32'd4231, -32'd7258, 32'd8077, 32'd5135},
{-32'd11854, -32'd6646, -32'd4110, 32'd4542},
{-32'd4826, 32'd3139, 32'd2360, -32'd55},
{-32'd1193, -32'd7440, -32'd10820, -32'd7208},
{32'd739, -32'd2552, 32'd4099, 32'd2041},
{32'd3198, 32'd1469, -32'd3942, 32'd4010},
{32'd4014, 32'd5525, 32'd5174, -32'd7386},
{-32'd6691, -32'd4832, -32'd7946, -32'd2641},
{-32'd6640, 32'd10391, 32'd2575, -32'd6842},
{32'd8705, 32'd3773, 32'd4210, -32'd1644},
{32'd5451, -32'd2697, -32'd4453, 32'd4873},
{32'd5551, 32'd7120, 32'd636, 32'd1617},
{32'd4430, 32'd4181, 32'd2829, 32'd236},
{-32'd9643, 32'd1808, 32'd5853, -32'd526},
{32'd1766, 32'd338, 32'd1192, -32'd11584},
{32'd3884, -32'd7952, -32'd7292, 32'd11708},
{-32'd1127, 32'd8357, 32'd7925, -32'd1740},
{32'd4420, 32'd7431, -32'd200, -32'd2046},
{-32'd7219, 32'd4248, 32'd800, 32'd11750},
{32'd959, -32'd8940, -32'd3853, 32'd3676},
{-32'd2891, 32'd1093, 32'd2894, -32'd1770},
{-32'd10486, -32'd5811, 32'd2072, -32'd9250},
{-32'd13078, 32'd4214, 32'd2382, -32'd2829},
{-32'd1006, 32'd10042, 32'd1409, -32'd176},
{-32'd12888, -32'd11460, -32'd9202, 32'd1247},
{32'd4107, 32'd11143, -32'd3119, -32'd288},
{32'd3640, -32'd6147, 32'd7276, 32'd2278},
{32'd2681, 32'd11116, 32'd908, -32'd7283},
{32'd8756, -32'd6662, -32'd4069, 32'd1373},
{32'd6428, -32'd533, 32'd3786, 32'd7464},
{32'd1734, -32'd265, -32'd1374, -32'd1147},
{32'd14877, 32'd451, -32'd4386, -32'd811},
{-32'd2031, 32'd1940, 32'd6499, -32'd922},
{32'd2710, 32'd849, -32'd793, -32'd3853},
{32'd2030, -32'd11478, -32'd1260, -32'd5728},
{32'd1144, -32'd1289, 32'd1818, -32'd1973},
{-32'd2396, 32'd2697, -32'd12308, -32'd770},
{-32'd17665, 32'd5380, -32'd6757, 32'd4027},
{-32'd1063, 32'd2742, -32'd2815, 32'd9542},
{-32'd1105, -32'd1969, -32'd8043, -32'd6917},
{32'd8239, -32'd2523, 32'd4304, -32'd4858},
{32'd486, -32'd1694, 32'd1801, -32'd6838},
{-32'd3316, -32'd10338, -32'd1762, -32'd2925},
{-32'd4693, -32'd316, 32'd4769, 32'd3901},
{-32'd6536, 32'd5034, -32'd12007, 32'd1422},
{32'd2750, 32'd2140, -32'd2561, -32'd946},
{-32'd4701, 32'd248, -32'd4716, 32'd1930},
{-32'd3501, -32'd10975, -32'd690, 32'd4698},
{32'd6385, -32'd1314, -32'd735, -32'd9727},
{-32'd9157, -32'd16080, -32'd6898, -32'd7396},
{-32'd11966, 32'd2392, 32'd4581, 32'd4321},
{32'd7747, 32'd4599, 32'd6038, -32'd352},
{32'd12467, -32'd2486, -32'd11313, 32'd3519},
{-32'd10509, -32'd550, 32'd2397, -32'd4982},
{-32'd497, -32'd3257, 32'd693, -32'd2084},
{32'd3290, -32'd9213, 32'd6657, 32'd5503},
{-32'd6323, 32'd393, 32'd3730, 32'd2710},
{32'd10127, -32'd11379, 32'd4064, -32'd2816},
{32'd5427, -32'd6776, 32'd7247, 32'd2133},
{32'd13362, 32'd7032, 32'd330, 32'd74},
{-32'd4074, -32'd2887, 32'd113, -32'd6419},
{-32'd9008, 32'd325, -32'd7901, 32'd5440},
{32'd926, -32'd4774, 32'd570, -32'd2637},
{32'd8215, 32'd71, 32'd2298, 32'd6747},
{32'd2047, -32'd7228, -32'd4416, -32'd4515},
{-32'd16934, -32'd7795, -32'd6473, 32'd640},
{32'd9537, 32'd8746, 32'd6015, -32'd2671},
{-32'd251, 32'd1915, -32'd413, -32'd1641},
{32'd16212, 32'd323, 32'd6899, -32'd674},
{32'd4971, 32'd863, -32'd5074, 32'd1148},
{-32'd817, -32'd11200, -32'd4800, -32'd7353},
{-32'd1677, 32'd5782, -32'd3479, 32'd690},
{-32'd7865, 32'd1824, 32'd1478, -32'd410},
{32'd1753, -32'd9674, 32'd3260, 32'd6699},
{-32'd2496, 32'd2922, -32'd4194, 32'd2956},
{32'd1579, -32'd475, -32'd1201, 32'd1152},
{-32'd4650, 32'd4822, -32'd653, 32'd631},
{32'd6978, 32'd13855, -32'd5270, 32'd1285},
{-32'd4021, 32'd3623, 32'd9404, 32'd1799},
{32'd11183, 32'd881, -32'd8957, 32'd7051},
{-32'd11903, 32'd3413, 32'd312, -32'd12833},
{32'd2981, -32'd6756, -32'd2374, -32'd5023},
{-32'd1693, 32'd2038, -32'd2826, 32'd2184},
{32'd6897, 32'd5639, 32'd8777, 32'd8681},
{32'd8588, 32'd11013, 32'd4380, -32'd4385},
{-32'd925, -32'd7598, -32'd4119, -32'd8964},
{-32'd16447, -32'd1518, -32'd2949, 32'd562},
{-32'd10614, -32'd8307, -32'd3306, 32'd4885},
{32'd1412, -32'd958, 32'd2992, -32'd2553},
{32'd16807, 32'd1875, -32'd4500, 32'd1749},
{-32'd2479, 32'd4642, -32'd3337, 32'd2155},
{32'd6482, 32'd17777, 32'd4661, -32'd5141},
{-32'd7879, -32'd2550, -32'd4323, -32'd7462},
{32'd12881, 32'd440, -32'd621, 32'd606},
{-32'd13070, 32'd7616, -32'd2525, 32'd2100},
{32'd8219, 32'd876, -32'd6543, 32'd11284},
{-32'd7236, -32'd13520, 32'd4556, -32'd4625},
{32'd11323, -32'd6106, -32'd1667, 32'd8543},
{32'd268, -32'd413, 32'd9600, -32'd3049},
{-32'd12138, -32'd463, -32'd3252, -32'd3728},
{-32'd313, -32'd5288, 32'd5973, 32'd1458},
{-32'd13311, 32'd7361, -32'd1374, -32'd6483},
{-32'd8380, 32'd1959, 32'd3956, -32'd5473},
{-32'd5920, 32'd1945, 32'd2308, -32'd2932},
{32'd487, 32'd7029, 32'd5794, 32'd34},
{32'd6474, 32'd2073, 32'd1379, 32'd2822},
{-32'd7475, 32'd1635, -32'd6770, -32'd2665}
},
{{32'd2945, 32'd742, 32'd9097, -32'd4816},
{32'd5594, 32'd14105, -32'd203, 32'd2120},
{32'd12514, 32'd8893, -32'd4801, 32'd5485},
{-32'd5471, 32'd14736, -32'd212, 32'd3555},
{-32'd686, -32'd2124, 32'd7982, -32'd1861},
{-32'd2391, -32'd8723, -32'd5353, 32'd6752},
{32'd1913, -32'd13647, 32'd2502, -32'd1814},
{-32'd4532, 32'd144, -32'd2247, -32'd12030},
{-32'd2503, -32'd4669, -32'd7776, -32'd5290},
{32'd4859, 32'd6226, 32'd3230, 32'd5318},
{-32'd4587, 32'd9213, 32'd11361, -32'd2533},
{-32'd332, 32'd1586, 32'd8021, 32'd3585},
{-32'd15820, 32'd6470, 32'd2131, -32'd4399},
{-32'd318, 32'd3502, 32'd37, -32'd336},
{-32'd3363, -32'd7823, -32'd4694, -32'd17484},
{32'd2505, 32'd7371, 32'd3959, -32'd13477},
{-32'd4091, 32'd6451, 32'd14722, 32'd3412},
{32'd1513, -32'd258, 32'd529, -32'd4632},
{-32'd4136, -32'd8253, -32'd7369, -32'd9642},
{-32'd15481, -32'd6395, -32'd898, 32'd3894},
{32'd5817, 32'd16627, -32'd6222, -32'd14607},
{-32'd6963, 32'd4545, -32'd10325, -32'd2249},
{32'd2520, -32'd4203, -32'd20751, -32'd4915},
{-32'd12165, -32'd4844, -32'd7129, 32'd5443},
{-32'd735, -32'd5225, -32'd6865, 32'd13095},
{-32'd3063, -32'd11831, 32'd4716, 32'd10},
{-32'd3526, -32'd6636, 32'd7075, -32'd6909},
{32'd4761, -32'd3877, -32'd10517, -32'd2062},
{-32'd8631, 32'd9873, 32'd5947, 32'd4349},
{-32'd926, -32'd8324, 32'd2130, -32'd4139},
{-32'd112, -32'd11639, -32'd4459, 32'd1110},
{-32'd16169, -32'd11769, 32'd1531, -32'd11021},
{32'd9282, -32'd1306, 32'd4766, -32'd3317},
{-32'd3913, 32'd11721, 32'd8479, -32'd1639},
{32'd1856, 32'd82, 32'd16573, 32'd8410},
{-32'd6274, -32'd8240, 32'd1431, 32'd1628},
{32'd12458, -32'd8871, -32'd10239, -32'd2366},
{-32'd10166, -32'd5657, 32'd8713, -32'd6283},
{-32'd11552, 32'd2198, 32'd7024, -32'd842},
{-32'd1255, 32'd11386, 32'd20735, 32'd12358},
{-32'd3955, 32'd15988, -32'd13157, -32'd3099},
{32'd2913, 32'd2501, 32'd725, 32'd5690},
{-32'd11852, 32'd5902, 32'd5467, -32'd4015},
{-32'd1112, 32'd1655, -32'd6839, -32'd1136},
{-32'd9867, -32'd164, 32'd10374, -32'd7003},
{32'd2867, 32'd5412, 32'd9324, 32'd1361},
{-32'd16296, -32'd2420, -32'd7607, -32'd5357},
{-32'd15745, -32'd3851, 32'd7481, -32'd4469},
{32'd677, -32'd5423, 32'd6752, 32'd9735},
{32'd8335, -32'd957, -32'd758, -32'd7882},
{-32'd4214, -32'd1760, 32'd3183, -32'd4464},
{-32'd3828, 32'd3079, 32'd9055, -32'd1894},
{32'd7278, 32'd1061, -32'd1055, 32'd772},
{-32'd2298, -32'd12829, -32'd1172, -32'd1771},
{32'd15568, -32'd15148, -32'd6397, -32'd137},
{32'd2600, 32'd9127, -32'd1085, 32'd2112},
{-32'd6260, -32'd2825, 32'd14239, 32'd7964},
{-32'd4457, -32'd8773, 32'd6452, -32'd4221},
{-32'd5284, 32'd2634, 32'd14408, -32'd2125},
{32'd7990, -32'd850, 32'd2575, 32'd1844},
{32'd10822, -32'd6783, -32'd9739, -32'd5372},
{-32'd6888, 32'd4230, 32'd15871, 32'd13472},
{-32'd4263, -32'd16214, 32'd2984, -32'd5980},
{32'd1275, 32'd4491, -32'd6113, -32'd1736},
{32'd11291, -32'd10877, -32'd7903, 32'd9010},
{-32'd5128, -32'd252, -32'd1808, 32'd4473},
{32'd6785, -32'd94, -32'd10525, -32'd7129},
{32'd3091, 32'd5502, 32'd5677, 32'd248},
{-32'd7147, -32'd1154, -32'd7271, -32'd11506},
{32'd15418, -32'd8814, 32'd5990, 32'd11457},
{32'd3349, 32'd2657, -32'd3413, 32'd2560},
{32'd5659, 32'd11625, 32'd5450, -32'd1432},
{-32'd3260, 32'd3176, -32'd2481, -32'd7168},
{-32'd9653, 32'd13234, -32'd3949, 32'd4292},
{32'd2897, -32'd2155, -32'd8038, -32'd628},
{32'd2831, 32'd5368, -32'd12595, 32'd465},
{32'd1179, -32'd2646, 32'd139, 32'd4333},
{32'd13524, -32'd4988, -32'd230, -32'd3174},
{32'd935, -32'd6344, 32'd2642, 32'd1073},
{32'd5678, -32'd7778, 32'd11482, 32'd7556},
{32'd6265, -32'd2212, 32'd6803, -32'd3067},
{32'd3724, -32'd3029, 32'd2710, 32'd3882},
{32'd2392, -32'd130, 32'd6365, -32'd5854},
{32'd14009, -32'd3705, -32'd1606, 32'd1445},
{32'd8849, -32'd5414, -32'd5761, 32'd2564},
{-32'd4767, -32'd11113, 32'd3895, -32'd7258},
{-32'd427, -32'd17098, 32'd13397, 32'd4579},
{-32'd9136, -32'd1460, 32'd782, -32'd5780},
{-32'd12345, 32'd1807, 32'd10500, 32'd529},
{32'd1413, 32'd5536, -32'd321, -32'd7865},
{-32'd3055, -32'd1106, 32'd11047, 32'd6673},
{32'd6611, -32'd1781, -32'd6848, -32'd4782},
{-32'd2317, -32'd532, -32'd4100, -32'd2527},
{32'd18021, -32'd977, 32'd3483, 32'd6701},
{-32'd6369, -32'd747, 32'd9293, -32'd15762},
{32'd6641, 32'd1411, -32'd7948, -32'd11807},
{32'd5570, 32'd6908, 32'd12283, 32'd2885},
{32'd10134, -32'd15415, -32'd12, -32'd7350},
{32'd5439, 32'd10505, -32'd11023, 32'd8438},
{32'd10307, 32'd4163, 32'd9943, -32'd4267},
{32'd1468, 32'd5718, -32'd4840, -32'd1253},
{-32'd4839, 32'd2261, 32'd101, -32'd10476},
{32'd4498, 32'd6827, 32'd20469, 32'd5893},
{32'd2757, 32'd6649, 32'd5888, 32'd14987},
{-32'd6193, 32'd9176, 32'd3603, 32'd427},
{32'd2275, 32'd525, 32'd6970, 32'd2533},
{-32'd3765, -32'd426, -32'd1627, -32'd375},
{-32'd3808, -32'd8945, -32'd728, -32'd2284},
{-32'd932, 32'd2407, 32'd2253, 32'd6004},
{-32'd4866, 32'd9836, 32'd17767, -32'd4465},
{32'd5896, 32'd5718, -32'd13542, 32'd7661},
{-32'd1470, 32'd10772, 32'd13098, 32'd4187},
{-32'd2735, -32'd8331, 32'd7863, 32'd10979},
{-32'd4109, -32'd4291, 32'd5337, 32'd0},
{32'd4851, -32'd8529, 32'd3995, -32'd16738},
{32'd8026, 32'd3763, -32'd26420, 32'd2566},
{-32'd10013, -32'd6795, 32'd3358, 32'd9000},
{32'd2762, -32'd10981, -32'd7980, -32'd28},
{32'd17837, 32'd7201, 32'd6679, -32'd11885},
{32'd6958, 32'd3403, 32'd2097, 32'd95},
{-32'd652, -32'd9880, -32'd3866, -32'd6801},
{32'd2364, 32'd1918, 32'd6469, 32'd5374},
{32'd10083, 32'd8053, -32'd9656, -32'd6993},
{-32'd2784, -32'd2073, -32'd8048, 32'd3277},
{-32'd1627, -32'd6885, 32'd510, -32'd3111},
{32'd12012, -32'd3671, 32'd4717, 32'd9042},
{-32'd3619, -32'd3500, 32'd2061, -32'd7681},
{-32'd8025, 32'd2210, -32'd5283, -32'd5116},
{-32'd1114, -32'd2154, 32'd3530, -32'd9554},
{-32'd4658, 32'd4259, 32'd2100, 32'd6129},
{-32'd14643, -32'd12000, -32'd3910, -32'd4928},
{-32'd6228, -32'd4334, 32'd11198, -32'd132},
{-32'd11211, -32'd2737, 32'd2611, 32'd7662},
{-32'd2779, 32'd2053, 32'd3371, -32'd1862},
{-32'd2607, 32'd12350, -32'd6270, -32'd13575},
{32'd11079, 32'd3704, -32'd7609, -32'd867},
{-32'd103, 32'd4913, -32'd13570, 32'd6234},
{32'd1635, 32'd5543, 32'd672, 32'd11159},
{32'd1174, -32'd1439, -32'd3398, -32'd3138},
{-32'd2023, -32'd11707, 32'd3718, -32'd3220},
{-32'd9112, -32'd3389, -32'd3281, 32'd1766},
{32'd11492, 32'd5881, -32'd892, 32'd6877},
{32'd4527, 32'd10787, -32'd4123, -32'd9709},
{32'd2998, -32'd8877, 32'd11563, -32'd8904},
{-32'd3709, -32'd6508, 32'd1100, 32'd12394},
{32'd15046, -32'd3611, 32'd4250, -32'd2611},
{-32'd1611, 32'd715, 32'd13009, 32'd801},
{-32'd11529, -32'd9517, -32'd1894, 32'd2711},
{32'd14074, 32'd9329, 32'd1891, 32'd1167},
{-32'd6026, -32'd8664, -32'd10811, -32'd5901},
{32'd3509, -32'd1698, 32'd1685, 32'd2196},
{32'd1647, -32'd7137, -32'd1782, 32'd3553},
{32'd7896, 32'd7512, -32'd7424, -32'd6193},
{32'd17686, 32'd4915, 32'd10264, -32'd6067},
{-32'd1640, 32'd5579, -32'd3343, 32'd1975},
{32'd6505, -32'd15745, 32'd491, -32'd11947},
{32'd589, 32'd6869, -32'd1211, -32'd823},
{-32'd8536, -32'd2110, 32'd11991, -32'd7251},
{-32'd508, 32'd3423, 32'd4229, -32'd6233},
{32'd2780, -32'd4325, 32'd8943, -32'd3755},
{32'd4898, -32'd6901, -32'd20529, -32'd9283},
{32'd6965, -32'd8608, -32'd14161, 32'd1660},
{-32'd1625, -32'd3145, -32'd2155, -32'd802},
{32'd2003, 32'd13061, 32'd3423, 32'd14303},
{32'd74, -32'd1274, 32'd8302, 32'd2187},
{32'd5862, -32'd5489, -32'd7038, 32'd341},
{32'd2065, -32'd12705, -32'd979, -32'd3383},
{-32'd6474, 32'd3949, 32'd2876, -32'd3454},
{-32'd3581, 32'd438, 32'd15274, -32'd888},
{-32'd2887, -32'd17206, -32'd8285, 32'd7094},
{-32'd7901, -32'd1289, 32'd2205, 32'd5175},
{-32'd0, 32'd13381, 32'd3686, 32'd3121},
{-32'd1868, 32'd9029, 32'd9722, 32'd6502},
{-32'd10837, -32'd8682, 32'd875, 32'd2098},
{32'd5102, -32'd1035, -32'd4606, -32'd4403},
{32'd5365, -32'd2400, 32'd6660, 32'd1249},
{-32'd8601, 32'd9095, 32'd14409, 32'd297},
{32'd3502, 32'd2249, -32'd11794, -32'd789},
{-32'd13008, -32'd1033, 32'd9014, -32'd1260},
{32'd1932, -32'd4027, -32'd6821, -32'd8967},
{-32'd17677, 32'd3355, -32'd2890, -32'd627},
{-32'd5496, -32'd4623, 32'd7385, -32'd1116},
{32'd14194, -32'd2973, -32'd16258, 32'd2034},
{32'd1847, 32'd10876, 32'd922, -32'd10376},
{32'd13014, -32'd1431, 32'd553, 32'd2273},
{32'd2852, 32'd2575, -32'd11895, -32'd4613},
{32'd759, 32'd6170, -32'd3358, 32'd3165},
{32'd10031, 32'd11157, 32'd3108, 32'd121},
{32'd6439, 32'd5689, -32'd8594, -32'd5470},
{-32'd308, -32'd1448, -32'd1792, -32'd3696},
{32'd5992, 32'd944, 32'd7120, 32'd3551},
{-32'd16440, -32'd2877, -32'd5188, -32'd2694},
{32'd6353, 32'd3246, 32'd6227, -32'd9830},
{-32'd6547, -32'd12243, 32'd6115, -32'd10791},
{32'd4172, 32'd3911, -32'd13475, -32'd3061},
{-32'd8835, 32'd1489, -32'd8720, 32'd12346},
{32'd8545, 32'd6986, 32'd6217, -32'd382},
{32'd19032, 32'd4506, -32'd7098, 32'd3744},
{32'd1117, -32'd549, 32'd3534, 32'd4259},
{-32'd1113, -32'd3506, 32'd2681, -32'd472},
{-32'd10119, -32'd2848, -32'd7228, -32'd2047},
{-32'd1098, 32'd4253, -32'd1696, -32'd12665},
{-32'd535, 32'd6950, -32'd2060, 32'd7562},
{32'd11545, -32'd1808, -32'd1599, -32'd8878},
{32'd5359, -32'd11020, -32'd1858, 32'd3977},
{-32'd6044, 32'd6146, 32'd13978, 32'd7420},
{32'd282, 32'd14935, -32'd5242, 32'd9148},
{32'd6214, -32'd6383, -32'd6634, -32'd12865},
{32'd594, -32'd7855, 32'd8596, 32'd3787},
{-32'd10323, 32'd3344, 32'd16184, -32'd2709},
{32'd8246, 32'd690, -32'd4296, 32'd5385},
{-32'd1718, -32'd15391, -32'd967, 32'd3688},
{32'd3071, -32'd10009, -32'd7767, 32'd1096},
{32'd5732, 32'd6112, -32'd8475, -32'd5474},
{32'd16855, 32'd3242, -32'd1591, -32'd5182},
{-32'd5558, -32'd7272, -32'd11225, 32'd509},
{32'd1131, -32'd1981, -32'd817, -32'd6477},
{-32'd409, -32'd4108, -32'd21101, -32'd11290},
{32'd10128, -32'd6118, 32'd12597, 32'd8833},
{32'd1210, -32'd692, -32'd10291, -32'd4702},
{32'd7555, 32'd2888, -32'd9893, 32'd6350},
{-32'd6156, 32'd2821, -32'd12103, -32'd432},
{32'd4975, 32'd577, 32'd3514, -32'd34},
{-32'd2362, -32'd12594, -32'd4586, -32'd7845},
{-32'd6866, 32'd5355, 32'd999, -32'd3419},
{32'd168, -32'd6330, 32'd8878, 32'd4445},
{32'd7134, 32'd10544, 32'd8725, -32'd8559},
{32'd6092, -32'd6652, -32'd7422, -32'd5348},
{-32'd10598, -32'd2362, 32'd12597, -32'd1542},
{-32'd10272, -32'd1810, -32'd8259, 32'd8222},
{-32'd14310, 32'd8891, 32'd1464, -32'd7218},
{-32'd4681, 32'd359, 32'd7312, -32'd11575},
{32'd6954, -32'd2694, -32'd5402, -32'd7235},
{32'd8105, -32'd10854, -32'd18637, 32'd2488},
{32'd11778, -32'd7470, -32'd7411, -32'd9968},
{32'd4947, -32'd5377, -32'd7156, -32'd9656},
{-32'd10289, 32'd3596, -32'd6206, -32'd7488},
{-32'd2815, 32'd8034, 32'd7252, -32'd6151},
{-32'd1598, 32'd10599, 32'd7528, 32'd5233},
{-32'd1231, 32'd1298, 32'd11402, -32'd3195},
{-32'd1166, 32'd1710, 32'd606, 32'd7278},
{32'd8946, -32'd4794, 32'd2205, -32'd1178},
{-32'd6149, -32'd11777, -32'd6993, -32'd393},
{32'd11418, 32'd5342, 32'd5101, 32'd5972},
{32'd9576, 32'd9695, 32'd7122, 32'd3712},
{32'd10995, 32'd9646, -32'd9262, -32'd3540},
{32'd3721, -32'd9053, 32'd112, -32'd12456},
{32'd2407, -32'd5913, -32'd15071, 32'd2134},
{32'd4072, 32'd273, -32'd3354, -32'd4780},
{32'd11219, -32'd4987, 32'd2480, 32'd98},
{32'd4314, 32'd1076, 32'd1501, -32'd5471},
{-32'd16360, -32'd8146, -32'd1392, -32'd6576},
{32'd7962, -32'd5708, 32'd193, 32'd7288},
{-32'd9655, -32'd1512, -32'd8114, -32'd4701},
{32'd814, -32'd7034, 32'd195, -32'd8522},
{32'd2812, -32'd4952, 32'd12593, 32'd9006},
{-32'd11659, 32'd13433, -32'd1252, 32'd9867},
{32'd3040, 32'd4403, -32'd4186, 32'd2175},
{-32'd19300, -32'd7841, 32'd7614, -32'd5676},
{32'd3413, -32'd471, 32'd4988, 32'd11168},
{-32'd11667, -32'd5476, 32'd3989, -32'd2237},
{-32'd5764, -32'd644, 32'd5083, -32'd240},
{32'd13880, -32'd9628, -32'd15734, 32'd19445},
{-32'd2457, 32'd351, 32'd1982, 32'd1090},
{-32'd3790, -32'd23, -32'd6020, -32'd8054},
{-32'd4816, -32'd6447, 32'd96, 32'd5929},
{32'd404, 32'd4253, 32'd4832, 32'd6832},
{32'd9173, -32'd5171, 32'd5307, -32'd596},
{-32'd9481, -32'd9062, 32'd1534, 32'd893},
{-32'd655, -32'd1217, -32'd11389, 32'd5255},
{32'd2064, -32'd2295, -32'd2744, 32'd1486},
{-32'd2559, -32'd1846, 32'd890, 32'd3886},
{-32'd8719, 32'd5663, 32'd3076, 32'd908},
{-32'd1787, -32'd553, -32'd7198, 32'd917},
{32'd1222, 32'd6052, -32'd184, -32'd586},
{32'd6055, -32'd1892, 32'd5081, 32'd8057},
{32'd4043, 32'd9236, 32'd7656, 32'd6675},
{-32'd9769, 32'd7054, 32'd1216, -32'd7908},
{32'd2934, -32'd4482, -32'd14746, -32'd4150},
{-32'd3049, 32'd6351, -32'd4184, -32'd3907},
{32'd8333, -32'd3210, -32'd5463, -32'd9920},
{32'd6174, 32'd5386, 32'd9720, -32'd5949},
{32'd3665, 32'd10372, 32'd14719, 32'd601},
{32'd11910, 32'd7129, -32'd10187, 32'd2052},
{32'd627, 32'd4485, -32'd3008, -32'd6803},
{32'd2445, -32'd5770, 32'd2860, -32'd1759},
{32'd8522, -32'd3504, -32'd5721, -32'd4743},
{32'd9607, -32'd19785, -32'd19424, -32'd9356},
{32'd1878, -32'd8371, -32'd16137, 32'd2323},
{-32'd8149, 32'd2253, -32'd3667, 32'd230},
{-32'd10514, -32'd5426, -32'd847, 32'd7414},
{32'd2928, 32'd7849, 32'd2556, 32'd9666},
{32'd4274, -32'd1229, 32'd10180, -32'd9454},
{-32'd9211, -32'd9171, -32'd2743, -32'd1671},
{-32'd3342, -32'd3179, 32'd680, 32'd16},
{32'd8644, -32'd5309, 32'd8827, -32'd6901},
{-32'd12500, -32'd530, 32'd7196, 32'd13610},
{-32'd872, 32'd7415, 32'd4887, -32'd848},
{32'd1602, 32'd9643, 32'd3802, 32'd1810},
{-32'd8799, -32'd1476, -32'd12054, -32'd12139}
},
{{-32'd6448, 32'd591, 32'd5570, 32'd4721},
{-32'd7640, 32'd13, -32'd970, -32'd2057},
{32'd2643, 32'd1243, 32'd1230, 32'd6328},
{32'd13019, 32'd2607, -32'd9544, 32'd5865},
{32'd7375, -32'd9129, -32'd4472, 32'd6073},
{32'd1450, -32'd6994, -32'd4238, 32'd2366},
{32'd4825, 32'd7115, 32'd601, 32'd10778},
{-32'd5130, -32'd7173, 32'd6260, -32'd1355},
{-32'd10950, -32'd1255, 32'd5041, -32'd6537},
{32'd7252, 32'd3871, 32'd1612, 32'd12001},
{32'd5281, 32'd3849, 32'd6844, -32'd630},
{-32'd825, -32'd7465, -32'd6119, -32'd3180},
{32'd5453, 32'd562, 32'd6403, 32'd136},
{32'd3671, 32'd12447, 32'd2944, 32'd782},
{-32'd3190, 32'd13484, 32'd255, 32'd1849},
{32'd6614, 32'd6915, 32'd7029, -32'd971},
{-32'd3764, -32'd1943, -32'd7430, 32'd6467},
{32'd2816, -32'd407, -32'd12624, -32'd3309},
{-32'd3842, -32'd3278, 32'd5348, 32'd220},
{-32'd3117, 32'd6725, -32'd523, 32'd2553},
{32'd7548, -32'd1137, 32'd3455, 32'd5156},
{-32'd437, -32'd583, -32'd1045, 32'd16},
{-32'd1472, 32'd9086, -32'd4193, -32'd56},
{32'd1713, 32'd3099, 32'd11948, -32'd2322},
{32'd7938, 32'd1556, 32'd1257, 32'd9501},
{32'd10609, -32'd100, -32'd1814, 32'd2071},
{-32'd8991, 32'd2093, 32'd469, 32'd1850},
{-32'd874, 32'd3350, -32'd6685, 32'd5139},
{32'd1845, -32'd1648, 32'd3891, 32'd3199},
{-32'd6960, -32'd18001, 32'd2927, -32'd4147},
{32'd7573, -32'd442, -32'd1964, -32'd1785},
{32'd2560, 32'd6246, 32'd3062, -32'd4850},
{32'd935, -32'd10407, 32'd5292, 32'd3023},
{-32'd1795, 32'd914, -32'd984, -32'd929},
{-32'd162, -32'd4189, -32'd936, 32'd4755},
{-32'd5686, 32'd15154, 32'd7484, -32'd1346},
{-32'd7083, -32'd4139, -32'd2756, 32'd9910},
{-32'd6776, 32'd4150, -32'd5166, 32'd5008},
{32'd12168, -32'd7707, -32'd561, 32'd6773},
{-32'd7043, -32'd14260, -32'd1881, -32'd2426},
{32'd4703, -32'd8411, -32'd5730, 32'd6548},
{-32'd1718, 32'd7102, 32'd12265, -32'd2388},
{32'd385, -32'd3074, -32'd8225, 32'd2886},
{32'd211, 32'd4991, 32'd3930, -32'd3559},
{-32'd12146, -32'd12894, 32'd1871, -32'd4414},
{-32'd14, -32'd16476, -32'd469, -32'd5891},
{-32'd667, 32'd3855, -32'd2691, -32'd1096},
{-32'd6630, -32'd8756, -32'd6839, -32'd3998},
{32'd8777, 32'd17251, 32'd847, -32'd2908},
{-32'd1400, -32'd4980, -32'd4256, -32'd2159},
{-32'd8470, -32'd2755, 32'd1064, 32'd6979},
{32'd4044, 32'd14771, -32'd472, -32'd3199},
{32'd6720, 32'd2139, 32'd2760, -32'd1043},
{32'd6352, -32'd979, 32'd4990, -32'd7197},
{-32'd124, -32'd1020, -32'd8769, -32'd2647},
{-32'd8355, 32'd5518, 32'd2086, -32'd3279},
{32'd9574, 32'd11713, -32'd6616, -32'd2389},
{32'd3106, -32'd1688, 32'd1411, -32'd3889},
{-32'd5816, -32'd15280, 32'd3172, -32'd4184},
{-32'd2568, 32'd2468, -32'd6378, -32'd5088},
{32'd5422, -32'd10450, -32'd8555, 32'd6020},
{32'd5112, 32'd2049, -32'd501, -32'd5418},
{-32'd13413, 32'd4118, 32'd4978, 32'd1600},
{32'd6800, 32'd1026, 32'd2787, 32'd901},
{-32'd3284, -32'd480, -32'd5813, 32'd2466},
{32'd350, -32'd1791, 32'd7552, 32'd8031},
{-32'd6332, -32'd8137, 32'd3066, 32'd4840},
{-32'd7423, 32'd650, 32'd694, -32'd7535},
{32'd2649, -32'd6619, 32'd394, 32'd4883},
{-32'd6480, -32'd3445, 32'd2047, -32'd1824},
{-32'd10365, -32'd751, -32'd4707, 32'd3632},
{-32'd2113, 32'd2338, 32'd4957, 32'd1303},
{-32'd768, 32'd4798, 32'd9539, -32'd2358},
{32'd9299, -32'd3732, -32'd6473, 32'd4870},
{32'd6846, -32'd5519, 32'd1762, 32'd2780},
{32'd6074, 32'd6945, 32'd8975, -32'd3910},
{32'd378, -32'd477, 32'd4285, -32'd315},
{-32'd257, -32'd9757, -32'd7173, 32'd13635},
{-32'd7144, 32'd5429, 32'd9558, 32'd4166},
{-32'd9151, -32'd173, -32'd1583, -32'd1007},
{32'd12399, -32'd3097, 32'd606, 32'd6645},
{32'd301, 32'd894, 32'd5248, 32'd4205},
{-32'd329, -32'd20587, 32'd494, -32'd886},
{32'd7467, 32'd3537, 32'd1624, 32'd5322},
{32'd3733, -32'd5589, 32'd3290, -32'd1287},
{-32'd2812, 32'd4655, 32'd5874, -32'd6320},
{32'd5107, 32'd582, -32'd8499, 32'd1888},
{32'd7463, -32'd2783, -32'd3154, -32'd4679},
{-32'd2891, -32'd6201, -32'd2492, -32'd927},
{-32'd9010, -32'd15573, -32'd5699, -32'd7611},
{32'd2635, 32'd8916, -32'd9328, -32'd203},
{32'd2072, -32'd241, 32'd5556, 32'd318},
{32'd10435, -32'd2208, 32'd1869, 32'd6312},
{32'd3608, 32'd2956, -32'd3390, 32'd6446},
{-32'd2947, -32'd7570, 32'd747, -32'd12940},
{-32'd6435, -32'd2697, 32'd6038, -32'd6785},
{32'd1644, -32'd8564, -32'd1124, 32'd6073},
{-32'd670, 32'd1795, 32'd5411, -32'd3951},
{32'd9555, -32'd566, 32'd3216, -32'd984},
{32'd8854, 32'd2510, 32'd2233, 32'd7928},
{-32'd321, -32'd4231, 32'd4910, -32'd6521},
{-32'd1328, -32'd2047, 32'd1219, -32'd298},
{-32'd11624, -32'd10811, 32'd5592, 32'd2642},
{-32'd2433, -32'd4175, -32'd4428, 32'd7007},
{32'd14276, -32'd4420, -32'd6806, -32'd1149},
{-32'd1478, -32'd3582, -32'd215, -32'd650},
{-32'd4305, 32'd5710, 32'd566, -32'd4128},
{32'd15130, -32'd3852, 32'd3449, 32'd6102},
{32'd4164, -32'd6696, 32'd10245, 32'd1892},
{32'd2197, 32'd5039, 32'd601, 32'd1232},
{32'd7360, 32'd1375, 32'd1104, 32'd9569},
{-32'd203, 32'd805, 32'd3072, 32'd2272},
{-32'd652, -32'd3158, 32'd2686, 32'd7847},
{32'd4944, 32'd13616, -32'd2619, 32'd2044},
{32'd4810, 32'd1514, 32'd7322, 32'd3565},
{32'd47, 32'd7576, 32'd1311, -32'd6228},
{32'd626, -32'd2026, -32'd7920, 32'd5610},
{-32'd5722, 32'd1768, 32'd1816, 32'd5460},
{32'd262, 32'd7734, 32'd2349, -32'd1051},
{32'd3800, 32'd13466, 32'd3190, 32'd6662},
{-32'd3084, 32'd6275, -32'd5316, 32'd2190},
{32'd9770, 32'd4354, 32'd5582, -32'd4632},
{-32'd2681, 32'd2187, -32'd6919, -32'd9077},
{-32'd6659, -32'd2759, -32'd5335, -32'd3674},
{32'd1573, -32'd13079, -32'd7558, -32'd3579},
{32'd2023, -32'd3237, 32'd9067, -32'd1031},
{-32'd9493, 32'd7757, -32'd5020, -32'd6324},
{-32'd6944, -32'd324, 32'd3564, 32'd1718},
{-32'd8595, 32'd816, 32'd0, -32'd712},
{-32'd2471, 32'd2807, -32'd6868, -32'd581},
{32'd6835, 32'd1698, -32'd5677, -32'd1311},
{-32'd6463, -32'd8892, 32'd843, -32'd3970},
{-32'd6475, -32'd5230, -32'd4544, -32'd3427},
{32'd6239, 32'd1777, 32'd6468, 32'd4644},
{-32'd7475, 32'd2601, -32'd2634, 32'd2501},
{-32'd7624, -32'd1293, -32'd5635, -32'd3507},
{-32'd12987, 32'd3326, 32'd13242, -32'd2706},
{32'd5471, 32'd1686, 32'd3519, -32'd2718},
{32'd10820, 32'd350, 32'd713, -32'd4471},
{-32'd8230, -32'd3574, -32'd1398, -32'd5526},
{32'd4664, 32'd15421, -32'd184, 32'd12649},
{-32'd4482, -32'd12327, 32'd4282, -32'd3571},
{-32'd4533, -32'd2493, 32'd2537, -32'd6227},
{32'd5209, 32'd1320, 32'd838, -32'd5249},
{-32'd5466, 32'd2825, -32'd673, 32'd4321},
{32'd4426, 32'd14128, -32'd2998, -32'd5803},
{-32'd8404, -32'd569, 32'd1291, -32'd5115},
{-32'd2263, -32'd10732, 32'd1366, -32'd6342},
{32'd1955, -32'd5196, 32'd3463, -32'd2940},
{-32'd1543, -32'd4114, -32'd6805, -32'd996},
{-32'd8688, 32'd807, 32'd5215, -32'd9135},
{-32'd3549, 32'd9827, 32'd2229, 32'd1591},
{-32'd4781, 32'd1743, -32'd1799, -32'd2406},
{32'd4352, -32'd9743, 32'd1332, 32'd5257},
{-32'd12671, -32'd7392, 32'd657, -32'd6081},
{32'd43, -32'd7113, -32'd2122, -32'd4569},
{32'd7903, -32'd1109, 32'd2300, 32'd1792},
{-32'd8571, -32'd2172, -32'd7605, -32'd10693},
{32'd2094, -32'd10005, -32'd8905, -32'd3778},
{-32'd3245, -32'd9854, 32'd14892, 32'd1462},
{-32'd6105, 32'd9280, 32'd809, 32'd634},
{-32'd1675, 32'd2141, 32'd4356, 32'd8427},
{-32'd10464, -32'd1725, -32'd1963, -32'd1548},
{-32'd1254, -32'd8710, -32'd6694, 32'd5100},
{-32'd20, 32'd166, -32'd1278, -32'd5931},
{-32'd3105, 32'd1537, 32'd3699, 32'd1616},
{-32'd1593, -32'd12767, 32'd1077, 32'd1386},
{-32'd3473, 32'd6893, 32'd125, -32'd4853},
{-32'd6997, -32'd8423, 32'd3186, -32'd7665},
{-32'd7278, 32'd12791, -32'd4884, -32'd9291},
{-32'd7276, 32'd782, 32'd4276, 32'd1262},
{32'd6569, -32'd1449, 32'd10581, -32'd5804},
{32'd3742, -32'd1936, -32'd4436, 32'd7429},
{32'd5488, -32'd5543, 32'd2563, 32'd145},
{-32'd1608, -32'd301, -32'd1456, 32'd7804},
{-32'd3267, 32'd712, 32'd12554, 32'd8985},
{-32'd9311, -32'd2249, -32'd5047, 32'd3277},
{32'd4433, -32'd6168, -32'd3631, 32'd1100},
{32'd1017, 32'd2124, 32'd1541, 32'd1549},
{32'd1093, -32'd11576, 32'd5070, -32'd3210},
{32'd2009, 32'd2124, 32'd2697, -32'd1700},
{-32'd401, -32'd4481, -32'd5832, -32'd2027},
{32'd8517, -32'd284, 32'd888, -32'd8853},
{-32'd16158, -32'd12345, -32'd821, 32'd296},
{-32'd6343, -32'd6215, -32'd4258, 32'd7482},
{32'd826, -32'd2165, -32'd5887, 32'd5606},
{-32'd1309, 32'd8379, 32'd2383, 32'd4390},
{32'd3490, 32'd4249, -32'd10275, -32'd5832},
{32'd12543, -32'd7912, -32'd32, -32'd2097},
{-32'd15570, -32'd4211, 32'd3896, -32'd11391},
{-32'd763, 32'd811, 32'd8832, -32'd7288},
{-32'd3744, 32'd7936, 32'd2796, 32'd4774},
{-32'd3194, -32'd9064, -32'd9718, -32'd10785},
{-32'd218, -32'd1146, 32'd4785, 32'd2439},
{-32'd1942, -32'd4525, -32'd2412, 32'd1848},
{32'd13020, 32'd904, -32'd5135, 32'd4044},
{32'd200, -32'd1985, -32'd2616, -32'd3603},
{-32'd3100, -32'd7423, 32'd6220, 32'd8762},
{-32'd779, -32'd3376, 32'd4936, 32'd2483},
{32'd244, 32'd2288, -32'd7281, -32'd1562},
{-32'd3773, 32'd573, 32'd1281, -32'd8767},
{32'd6857, -32'd365, -32'd6747, 32'd1608},
{32'd10178, 32'd2501, 32'd1739, 32'd5945},
{32'd8540, 32'd12476, -32'd1156, 32'd7684},
{32'd4838, -32'd3893, 32'd4024, -32'd3004},
{-32'd8555, -32'd7370, -32'd6215, 32'd4798},
{32'd2924, 32'd626, 32'd921, 32'd11850},
{32'd4524, -32'd5210, -32'd136, 32'd1257},
{32'd2763, 32'd5181, -32'd16647, 32'd3923},
{32'd1103, -32'd16252, -32'd3587, -32'd7938},
{32'd4010, 32'd13335, 32'd1354, -32'd2089},
{-32'd1908, 32'd4923, -32'd7572, 32'd394},
{-32'd7424, 32'd7896, 32'd5836, -32'd545},
{32'd5096, -32'd3257, -32'd6663, 32'd611},
{32'd6413, -32'd2071, 32'd225, 32'd5293},
{-32'd7804, -32'd2298, -32'd4244, -32'd2718},
{32'd2891, -32'd5014, 32'd5364, 32'd1322},
{-32'd1656, -32'd5703, -32'd1646, 32'd1302},
{-32'd8672, -32'd4473, 32'd1712, -32'd1750},
{-32'd3011, 32'd564, 32'd7860, 32'd2233},
{-32'd4474, 32'd1850, -32'd4140, -32'd3435},
{-32'd3053, 32'd6717, -32'd961, 32'd10069},
{32'd3374, -32'd5481, -32'd287, 32'd5340},
{-32'd6902, 32'd4508, -32'd7713, 32'd1068},
{32'd1729, -32'd1844, -32'd841, -32'd2084},
{32'd8274, -32'd13569, 32'd3712, 32'd1332},
{-32'd4807, -32'd3789, -32'd2333, -32'd6768},
{-32'd1857, 32'd2398, 32'd7145, 32'd1791},
{-32'd6845, 32'd8474, -32'd42, 32'd1897},
{-32'd1997, 32'd2430, -32'd3515, -32'd821},
{-32'd7211, 32'd13923, -32'd939, -32'd776},
{-32'd10417, 32'd8107, -32'd9007, 32'd2729},
{32'd8096, 32'd10203, 32'd4358, 32'd264},
{32'd14540, 32'd3510, -32'd1514, 32'd6489},
{-32'd2608, -32'd5253, 32'd2231, -32'd4282},
{-32'd2056, 32'd10365, 32'd57, -32'd2937},
{-32'd15230, 32'd8836, -32'd6463, 32'd7129},
{32'd5123, -32'd7382, -32'd4157, -32'd5666},
{32'd778, -32'd6632, -32'd3470, -32'd61},
{-32'd4307, 32'd4186, 32'd15682, -32'd4115},
{-32'd125, 32'd11355, 32'd7595, -32'd9057},
{-32'd1091, 32'd2818, 32'd2963, -32'd4768},
{-32'd2494, -32'd8624, -32'd3585, -32'd5066},
{32'd4533, 32'd5244, 32'd7737, 32'd5549},
{32'd6719, 32'd2033, -32'd435, 32'd7442},
{32'd3772, -32'd6851, 32'd2152, -32'd6170},
{-32'd5541, -32'd9121, 32'd6029, -32'd7250},
{-32'd1518, -32'd11800, -32'd5712, -32'd4857},
{-32'd5639, -32'd8693, 32'd338, -32'd3720},
{32'd2861, -32'd10431, -32'd2600, 32'd2491},
{-32'd15721, 32'd9108, 32'd8615, -32'd909},
{-32'd4409, 32'd715, -32'd10252, 32'd1093},
{32'd759, -32'd4695, -32'd4507, -32'd3529},
{32'd614, 32'd7641, 32'd1092, 32'd9763},
{-32'd210, -32'd1578, -32'd981, -32'd4622},
{-32'd12648, 32'd5014, -32'd1600, 32'd1661},
{32'd3828, -32'd6967, 32'd8616, -32'd2109},
{32'd5583, 32'd7422, -32'd875, 32'd4675},
{-32'd15310, -32'd2846, -32'd7069, -32'd4472},
{32'd1932, -32'd1872, 32'd4063, 32'd797},
{32'd2256, 32'd1311, -32'd2980, -32'd1050},
{32'd316, -32'd2777, -32'd3110, -32'd438},
{32'd2380, 32'd11423, -32'd7213, -32'd662},
{32'd12843, -32'd7176, 32'd1314, -32'd4139},
{32'd8518, 32'd13710, -32'd4753, 32'd5121},
{32'd5205, -32'd4103, -32'd2106, -32'd2953},
{32'd6915, 32'd163, -32'd1034, -32'd514},
{-32'd53, 32'd3552, 32'd2791, 32'd952},
{-32'd7172, 32'd1247, 32'd1766, -32'd4700},
{32'd9316, -32'd764, 32'd1870, -32'd2366},
{-32'd2908, -32'd16832, -32'd187, 32'd3916},
{32'd3981, 32'd767, -32'd3480, 32'd3412},
{-32'd642, -32'd8203, -32'd12650, -32'd1567},
{-32'd4347, 32'd4004, 32'd3075, -32'd5114},
{32'd2961, -32'd3067, -32'd3536, -32'd4882},
{32'd7410, -32'd5894, 32'd1343, 32'd5266},
{32'd6801, 32'd5054, 32'd2396, 32'd10940},
{32'd9644, -32'd3906, -32'd2085, -32'd4383},
{32'd421, -32'd10019, -32'd5118, -32'd8028},
{-32'd991, -32'd3914, -32'd4817, -32'd3932},
{32'd3572, 32'd1094, 32'd911, 32'd4034},
{-32'd8611, 32'd7255, 32'd6115, -32'd565},
{32'd3245, 32'd6151, -32'd4426, 32'd3328},
{-32'd6146, 32'd1500, 32'd6279, 32'd8957},
{-32'd2825, 32'd402, -32'd6526, 32'd6413},
{-32'd1836, -32'd2454, 32'd7664, -32'd3487},
{32'd3064, 32'd3598, 32'd4788, 32'd2959},
{32'd9174, 32'd3919, 32'd10129, -32'd1447},
{32'd13200, 32'd10593, 32'd7375, -32'd3840},
{32'd4333, 32'd789, 32'd2221, -32'd5990},
{32'd12150, -32'd2073, -32'd1480, 32'd5235},
{32'd10882, 32'd11521, -32'd1059, 32'd9453},
{32'd4462, 32'd11739, 32'd3715, 32'd8475},
{32'd1819, 32'd3134, -32'd273, -32'd1254},
{-32'd9447, 32'd7506, -32'd1275, -32'd4994},
{-32'd8146, -32'd359, -32'd2804, -32'd10227},
{-32'd737, -32'd5669, -32'd3421, -32'd9313},
{32'd2017, -32'd8732, 32'd9185, 32'd3894},
{32'd6726, -32'd3187, -32'd4219, 32'd10119},
{32'd5372, 32'd15172, -32'd3867, 32'd5559}
},
{{32'd6349, 32'd4934, 32'd3281, 32'd1451},
{-32'd547, -32'd6829, -32'd12246, 32'd2591},
{-32'd1821, 32'd5384, -32'd2324, -32'd2265},
{32'd13548, 32'd4959, -32'd623, 32'd1902},
{-32'd9948, -32'd1689, -32'd7651, -32'd5293},
{32'd2002, -32'd2936, 32'd8861, 32'd3488},
{32'd20261, -32'd267, -32'd4664, -32'd6095},
{32'd3818, -32'd8973, -32'd7931, 32'd4203},
{-32'd6680, -32'd6291, 32'd255, -32'd1255},
{32'd2824, 32'd7008, 32'd13616, 32'd2160},
{-32'd6893, -32'd2490, -32'd3359, -32'd7320},
{32'd392, 32'd12817, 32'd8185, -32'd1103},
{-32'd333, -32'd11935, 32'd607, 32'd2751},
{32'd9602, 32'd2541, -32'd9717, -32'd2341},
{-32'd2986, 32'd463, -32'd6118, -32'd4383},
{-32'd5302, -32'd8542, -32'd1478, -32'd6862},
{32'd13338, -32'd4094, 32'd4221, 32'd389},
{-32'd5889, 32'd1652, -32'd2503, -32'd7965},
{-32'd7098, -32'd7320, 32'd1937, 32'd3421},
{32'd1506, 32'd4466, 32'd6698, 32'd791},
{-32'd5378, -32'd6428, -32'd37, 32'd1591},
{-32'd4575, 32'd753, -32'd3178, 32'd3185},
{-32'd6451, -32'd6564, 32'd1060, -32'd2814},
{-32'd11821, -32'd13616, -32'd7141, -32'd2373},
{32'd4475, -32'd1148, 32'd10434, -32'd1231},
{32'd15730, 32'd12148, -32'd5753, -32'd6118},
{-32'd1914, 32'd6012, -32'd2234, 32'd3503},
{-32'd13973, -32'd6272, -32'd3945, 32'd2995},
{32'd9831, 32'd11193, 32'd11710, -32'd3234},
{32'd2356, -32'd5573, -32'd5982, 32'd1739},
{-32'd18702, 32'd4417, -32'd9342, -32'd2193},
{-32'd3355, 32'd534, -32'd9696, -32'd9454},
{32'd956, 32'd15347, -32'd1215, 32'd2305},
{-32'd8814, -32'd6136, -32'd7999, -32'd276},
{-32'd6446, 32'd7479, 32'd8662, 32'd2345},
{32'd5105, -32'd443, 32'd1175, 32'd3387},
{-32'd169, 32'd4201, -32'd3466, -32'd2333},
{32'd7405, -32'd4884, 32'd2707, -32'd177},
{32'd6999, -32'd14714, 32'd465, -32'd6351},
{-32'd12538, -32'd4498, 32'd2827, -32'd930},
{-32'd5187, -32'd9661, 32'd4733, -32'd1166},
{-32'd4135, -32'd4643, -32'd7502, -32'd3828},
{-32'd8039, -32'd5155, -32'd5085, -32'd1668},
{-32'd8953, -32'd21121, -32'd17153, 32'd1301},
{-32'd11276, -32'd3967, -32'd2794, 32'd2355},
{-32'd6569, -32'd5853, -32'd11786, -32'd144},
{-32'd198, 32'd10101, -32'd4379, 32'd3081},
{32'd6733, -32'd1445, -32'd9598, 32'd1289},
{32'd16706, 32'd1316, 32'd1480, -32'd966},
{32'd4560, 32'd4164, -32'd3318, -32'd558},
{32'd2917, 32'd162, 32'd4160, -32'd4073},
{32'd4057, 32'd6189, 32'd478, -32'd509},
{32'd7867, 32'd14491, -32'd7107, -32'd9630},
{-32'd6807, -32'd6362, 32'd6508, 32'd1662},
{-32'd4528, -32'd4856, -32'd4119, -32'd4582},
{-32'd13313, -32'd4994, -32'd1953, 32'd3365},
{32'd11535, 32'd7089, 32'd3300, 32'd1345},
{32'd2751, -32'd9588, -32'd5064, -32'd8182},
{-32'd1886, -32'd4843, -32'd1377, -32'd422},
{-32'd1521, 32'd2787, -32'd3137, 32'd2530},
{-32'd4271, -32'd1443, -32'd5007, 32'd490},
{-32'd704, -32'd1475, 32'd6222, 32'd3087},
{-32'd6527, -32'd11037, -32'd12892, -32'd2809},
{32'd6321, 32'd2800, -32'd2724, 32'd6241},
{-32'd2244, 32'd4558, -32'd2329, 32'd4648},
{32'd1493, 32'd4127, 32'd5723, -32'd1064},
{32'd3538, -32'd3439, 32'd5298, 32'd1462},
{-32'd7645, 32'd6819, -32'd11861, -32'd2334},
{32'd2589, -32'd13108, -32'd49, -32'd1017},
{32'd7848, -32'd2895, 32'd2474, 32'd7654},
{32'd4381, 32'd26, -32'd5478, -32'd1717},
{32'd797, -32'd10550, 32'd10774, -32'd2541},
{-32'd7035, -32'd1502, -32'd4171, -32'd3923},
{-32'd5607, -32'd11707, -32'd12144, -32'd502},
{32'd11344, 32'd3759, -32'd303, 32'd414},
{32'd8227, -32'd5935, -32'd574, 32'd9122},
{-32'd13372, -32'd5550, -32'd7873, 32'd3300},
{32'd7188, -32'd5854, -32'd6991, -32'd9358},
{32'd1484, -32'd2170, -32'd2411, 32'd1948},
{-32'd3493, -32'd990, -32'd3307, -32'd4504},
{-32'd6993, 32'd2113, 32'd7118, 32'd1728},
{-32'd7760, -32'd496, 32'd3173, 32'd3775},
{-32'd2952, -32'd6656, -32'd1308, -32'd3270},
{-32'd3441, 32'd2334, 32'd8643, -32'd6891},
{-32'd15813, -32'd2880, -32'd4317, -32'd3169},
{-32'd9017, -32'd14040, 32'd4110, -32'd2441},
{32'd2004, 32'd6645, 32'd7188, -32'd7141},
{-32'd13580, -32'd14013, -32'd1290, -32'd2456},
{32'd6865, -32'd3126, -32'd3245, -32'd737},
{-32'd10881, 32'd7777, -32'd7380, -32'd3249},
{32'd4735, 32'd70, 32'd11553, 32'd3978},
{-32'd10957, -32'd11597, -32'd12183, -32'd6088},
{-32'd11119, 32'd1785, 32'd6695, 32'd2528},
{32'd9467, 32'd10912, 32'd2874, -32'd3307},
{32'd7911, -32'd713, -32'd1912, -32'd5554},
{32'd2507, -32'd555, -32'd11468, -32'd276},
{32'd601, 32'd3233, 32'd10276, 32'd2984},
{-32'd7753, -32'd2402, 32'd1148, -32'd3391},
{-32'd6627, 32'd2808, -32'd1792, 32'd1007},
{32'd8950, 32'd7901, 32'd2626, -32'd323},
{-32'd6416, 32'd14578, -32'd6826, -32'd439},
{-32'd11351, 32'd2432, -32'd5083, -32'd2806},
{32'd2213, 32'd12666, -32'd1801, 32'd969},
{-32'd10328, 32'd5919, 32'd3873, -32'd3085},
{-32'd7208, -32'd10913, 32'd4967, -32'd895},
{32'd2038, 32'd2560, -32'd7795, -32'd1692},
{-32'd3986, 32'd768, -32'd1541, -32'd756},
{-32'd20059, -32'd4104, 32'd1129, -32'd2812},
{-32'd8360, -32'd883, -32'd3174, -32'd635},
{32'd793, 32'd309, -32'd5071, -32'd167},
{-32'd8905, -32'd10910, -32'd3418, -32'd507},
{32'd940, -32'd4955, 32'd5843, 32'd2662},
{-32'd71, -32'd11697, 32'd2443, 32'd6275},
{-32'd3844, 32'd2408, -32'd5904, 32'd264},
{-32'd6770, 32'd5627, -32'd2359, -32'd8909},
{32'd2188, 32'd2824, 32'd1721, 32'd3204},
{32'd6838, 32'd843, 32'd7062, -32'd1427},
{-32'd6484, 32'd6426, -32'd4996, 32'd7559},
{32'd2393, -32'd2918, -32'd1702, 32'd8072},
{32'd3045, 32'd18547, 32'd5715, 32'd5883},
{32'd5482, -32'd2514, -32'd3089, -32'd2223},
{32'd2783, -32'd962, -32'd10745, 32'd403},
{32'd369, 32'd1534, 32'd454, 32'd800},
{32'd20508, 32'd4167, 32'd1636, -32'd4497},
{32'd1118, -32'd1441, -32'd697, 32'd125},
{-32'd349, 32'd5461, -32'd6189, 32'd874},
{32'd2126, -32'd12303, -32'd2193, -32'd2947},
{-32'd17544, -32'd3571, 32'd1596, -32'd5447},
{-32'd447, 32'd673, -32'd12779, -32'd627},
{32'd9310, -32'd10681, -32'd652, 32'd2620},
{-32'd11791, 32'd5196, 32'd3484, -32'd990},
{-32'd7365, -32'd4132, -32'd4183, -32'd116},
{-32'd180, -32'd7645, -32'd1930, 32'd1831},
{32'd1989, 32'd13891, -32'd2497, -32'd1291},
{32'd968, 32'd5378, 32'd10276, 32'd5557},
{32'd3289, -32'd3845, 32'd7163, 32'd341},
{-32'd7586, 32'd401, 32'd3197, 32'd4759},
{-32'd9436, 32'd12037, 32'd2893, 32'd3382},
{-32'd7030, -32'd7211, -32'd5437, 32'd4035},
{32'd6948, -32'd5026, -32'd13675, -32'd2643},
{-32'd4123, -32'd6153, 32'd2244, -32'd493},
{-32'd6467, -32'd2222, -32'd10683, -32'd3460},
{32'd20010, 32'd4248, 32'd389, 32'd850},
{-32'd9192, 32'd3897, -32'd3565, -32'd7124},
{-32'd9093, 32'd9577, 32'd2946, 32'd2019},
{-32'd7747, -32'd3048, -32'd544, 32'd1011},
{-32'd25033, -32'd4679, -32'd13440, 32'd3151},
{-32'd12434, -32'd4313, 32'd3400, 32'd7248},
{32'd12423, 32'd11899, 32'd5611, 32'd6848},
{-32'd8716, -32'd7424, -32'd4785, 32'd6616},
{-32'd3373, -32'd8990, -32'd12034, 32'd3253},
{-32'd4590, 32'd446, 32'd1685, 32'd9488},
{-32'd18178, 32'd4210, -32'd305, -32'd2339},
{32'd9286, 32'd8784, -32'd3565, 32'd1139},
{-32'd3908, -32'd9617, -32'd8002, 32'd989},
{32'd12277, 32'd7496, 32'd4119, -32'd586},
{-32'd10374, 32'd595, 32'd7918, -32'd3494},
{32'd7032, -32'd8658, 32'd10724, 32'd803},
{-32'd23440, -32'd8198, 32'd4083, 32'd4556},
{-32'd3767, -32'd3727, 32'd9823, 32'd6239},
{32'd169, 32'd2955, -32'd6793, -32'd4865},
{32'd11327, 32'd5581, 32'd3968, 32'd1265},
{-32'd7551, -32'd1700, 32'd4542, -32'd1227},
{32'd9579, -32'd569, 32'd3683, 32'd1806},
{-32'd8256, -32'd2181, 32'd2842, -32'd222},
{32'd6365, 32'd1236, -32'd614, -32'd399},
{-32'd4245, 32'd5784, -32'd7013, -32'd8314},
{-32'd10986, -32'd1778, 32'd4816, 32'd475},
{32'd2735, 32'd11424, 32'd2672, 32'd1598},
{32'd10274, -32'd5264, -32'd9050, -32'd3305},
{-32'd800, -32'd15042, -32'd3420, -32'd4427},
{32'd9736, 32'd11320, -32'd9206, 32'd1466},
{32'd2540, 32'd18776, 32'd10247, 32'd5395},
{32'd18955, 32'd7842, -32'd4259, -32'd8966},
{32'd1953, -32'd4844, -32'd2154, 32'd8176},
{-32'd6751, -32'd11088, -32'd1671, 32'd7696},
{32'd943, 32'd1195, -32'd2921, 32'd8842},
{-32'd6713, -32'd4794, 32'd9145, 32'd8411},
{-32'd8173, 32'd441, -32'd5194, 32'd5659},
{32'd12676, -32'd2518, -32'd7132, -32'd3777},
{-32'd16988, -32'd1056, 32'd6779, 32'd263},
{-32'd9582, -32'd3740, 32'd3971, 32'd1086},
{32'd2066, 32'd5075, -32'd984, -32'd1730},
{-32'd649, -32'd10243, 32'd2445, -32'd955},
{-32'd10338, 32'd8751, 32'd3834, -32'd4937},
{32'd15429, -32'd7257, 32'd3157, 32'd990},
{32'd13057, 32'd5022, 32'd7843, 32'd2974},
{32'd2383, 32'd2026, 32'd1807, 32'd955},
{-32'd6122, -32'd8451, 32'd11799, 32'd263},
{-32'd3089, -32'd5030, 32'd3765, -32'd2642},
{32'd4652, -32'd2868, 32'd5341, 32'd8404},
{-32'd1767, -32'd10715, -32'd4952, -32'd5702},
{-32'd4653, -32'd5054, 32'd2800, -32'd6209},
{-32'd13027, 32'd2912, -32'd5442, -32'd4695},
{-32'd15259, 32'd7084, -32'd5637, -32'd2376},
{-32'd10000, 32'd6069, -32'd7923, 32'd1225},
{32'd9185, -32'd853, -32'd10648, 32'd811},
{-32'd14240, -32'd6108, 32'd4713, -32'd5573},
{-32'd6138, -32'd4007, 32'd2100, 32'd2717},
{32'd5070, 32'd6792, 32'd13633, -32'd698},
{32'd7070, -32'd2216, -32'd4495, 32'd1332},
{32'd2966, -32'd505, -32'd229, -32'd778},
{32'd5648, -32'd2888, 32'd9024, 32'd9271},
{32'd1740, 32'd9217, -32'd229, 32'd4408},
{-32'd7381, -32'd5099, 32'd1399, 32'd827},
{-32'd11745, 32'd8560, 32'd5997, -32'd1402},
{32'd4405, 32'd6154, 32'd8628, -32'd1384},
{-32'd17641, -32'd13124, 32'd530, -32'd373},
{32'd1675, -32'd382, 32'd3280, 32'd1785},
{-32'd8743, 32'd6326, 32'd6756, 32'd1578},
{-32'd23875, 32'd1147, -32'd301, -32'd1486},
{32'd95, -32'd4800, 32'd3977, 32'd300},
{-32'd13909, -32'd6264, -32'd234, -32'd3858},
{32'd7279, -32'd5004, -32'd21, 32'd327},
{32'd14184, 32'd6678, -32'd8057, -32'd583},
{32'd3623, -32'd3918, -32'd1816, -32'd3119},
{-32'd5113, 32'd4, 32'd5798, 32'd5657},
{-32'd2113, -32'd12005, -32'd9025, -32'd1065},
{32'd5115, 32'd2349, -32'd1284, 32'd11026},
{-32'd10456, 32'd874, -32'd2128, -32'd1506},
{32'd4754, -32'd5538, -32'd2889, -32'd1749},
{-32'd6819, -32'd862, 32'd7729, -32'd1781},
{-32'd7071, 32'd4785, -32'd1438, -32'd249},
{32'd3613, 32'd6517, 32'd884, 32'd1244},
{-32'd8271, -32'd344, 32'd4243, 32'd105},
{-32'd14968, 32'd597, 32'd1386, 32'd7084},
{32'd538, 32'd104, -32'd3281, -32'd2481},
{32'd10062, -32'd8267, -32'd5936, -32'd3820},
{32'd8604, -32'd1087, -32'd2956, -32'd8633},
{32'd8347, 32'd13157, 32'd8891, 32'd1059},
{-32'd13367, 32'd5582, -32'd1204, -32'd43},
{32'd5948, -32'd9652, -32'd7524, -32'd5314},
{32'd12543, 32'd857, -32'd1682, 32'd663},
{-32'd9337, 32'd2505, 32'd11032, -32'd3907},
{-32'd12372, -32'd7298, -32'd13480, 32'd7307},
{-32'd2814, 32'd995, -32'd9663, 32'd2643},
{-32'd2548, 32'd275, 32'd1077, -32'd9012},
{-32'd8200, 32'd10908, -32'd7850, -32'd3113},
{32'd5625, 32'd12530, -32'd4835, 32'd6889},
{-32'd9926, -32'd15206, -32'd1473, -32'd1548},
{-32'd1423, -32'd4375, 32'd331, -32'd5255},
{-32'd4593, 32'd3676, -32'd9298, 32'd2012},
{-32'd4131, -32'd11454, -32'd13073, -32'd4643},
{32'd5232, 32'd2679, 32'd1716, -32'd3615},
{-32'd1486, 32'd4394, 32'd10014, 32'd6722},
{32'd1165, 32'd6836, -32'd6882, 32'd7422},
{-32'd8358, -32'd5129, -32'd11630, -32'd7282},
{-32'd12262, 32'd3706, 32'd3964, -32'd3340},
{32'd163, 32'd14340, -32'd1552, 32'd1173},
{-32'd5402, 32'd2852, -32'd850, 32'd1623},
{-32'd7395, -32'd8412, -32'd4911, -32'd5111},
{-32'd7917, 32'd6546, 32'd4089, -32'd4745},
{32'd10192, -32'd2637, 32'd3794, 32'd2000},
{32'd73, -32'd1232, -32'd8331, -32'd1839},
{32'd2434, -32'd1642, -32'd2126, -32'd3726},
{32'd13702, 32'd6256, 32'd5788, 32'd445},
{-32'd5384, -32'd3767, -32'd53, 32'd4222},
{32'd15713, 32'd211, 32'd3948, 32'd10700},
{32'd2814, -32'd10685, -32'd3357, -32'd5393},
{32'd6659, 32'd9919, -32'd4080, 32'd3179},
{32'd12470, 32'd3368, 32'd11009, 32'd2633},
{-32'd8668, -32'd15262, 32'd5692, -32'd630},
{-32'd3453, -32'd232, -32'd6218, -32'd2547},
{32'd611, 32'd6464, -32'd1541, -32'd11778},
{-32'd6005, -32'd3378, -32'd2591, 32'd1137},
{32'd1968, 32'd1618, 32'd9353, 32'd1126},
{32'd19801, -32'd1607, -32'd2822, -32'd1481},
{-32'd9442, -32'd2303, 32'd5216, -32'd4298},
{32'd8503, -32'd6722, -32'd5704, -32'd4056},
{-32'd1602, 32'd9079, 32'd4992, -32'd7366},
{-32'd9369, -32'd5235, -32'd423, 32'd6555},
{32'd167, -32'd7108, 32'd2363, 32'd288},
{-32'd8253, -32'd7116, -32'd5304, 32'd4502},
{-32'd17310, -32'd692, -32'd4785, -32'd1963},
{32'd4072, 32'd5846, -32'd6105, -32'd1372},
{-32'd1730, -32'd2205, -32'd7815, -32'd5892},
{32'd2203, 32'd7814, 32'd13949, 32'd2170},
{-32'd5368, 32'd1667, -32'd142, 32'd149},
{-32'd6099, -32'd13080, -32'd12129, -32'd692},
{32'd3790, 32'd2666, 32'd4981, -32'd2810},
{32'd2425, -32'd1659, 32'd8935, 32'd1081},
{32'd5462, -32'd1349, -32'd2066, 32'd1424},
{32'd10648, 32'd5299, -32'd6616, -32'd3624},
{32'd1118, 32'd900, -32'd665, -32'd2553},
{-32'd1210, 32'd2307, 32'd15457, 32'd1278},
{32'd15694, 32'd3769, 32'd1103, -32'd2521},
{32'd12976, -32'd8181, -32'd2253, 32'd5006},
{-32'd12750, 32'd5359, 32'd1233, -32'd4981},
{32'd167, -32'd10644, -32'd2269, 32'd214},
{-32'd17419, -32'd20172, -32'd4891, 32'd5413},
{-32'd22032, 32'd450, 32'd4595, -32'd1180},
{32'd6759, 32'd10014, 32'd11695, 32'd3151},
{32'd7117, -32'd5197, 32'd82, -32'd4286},
{-32'd11201, -32'd11421, 32'd1287, 32'd2185},
{32'd5832, -32'd4803, 32'd5690, -32'd703},
{-32'd4693, -32'd5551, -32'd8138, -32'd2445},
{-32'd3864, 32'd1793, -32'd7210, -32'd1189},
{32'd598, 32'd1551, 32'd13761, 32'd8336},
{32'd197, 32'd6890, 32'd438, -32'd4260},
{32'd2589, -32'd14350, -32'd3755, 32'd7507}
},
{{32'd1865, 32'd13221, 32'd9510, 32'd5779},
{-32'd5275, -32'd7448, -32'd8729, 32'd971},
{32'd3086, 32'd3295, 32'd2834, 32'd2616},
{-32'd3611, 32'd5112, -32'd2045, 32'd2772},
{32'd11907, 32'd14352, -32'd5679, 32'd5281},
{-32'd9988, -32'd2082, 32'd10000, -32'd9443},
{32'd9592, 32'd3770, -32'd118, 32'd6227},
{-32'd4678, -32'd3097, -32'd33, 32'd4877},
{32'd265, 32'd5613, -32'd2011, -32'd609},
{32'd7616, 32'd12762, 32'd5143, 32'd112},
{-32'd1661, -32'd13715, 32'd12008, 32'd802},
{-32'd4121, 32'd4390, -32'd6915, 32'd6794},
{-32'd4024, 32'd1981, -32'd6884, -32'd1434},
{32'd8580, -32'd1683, -32'd11529, 32'd1227},
{32'd1748, -32'd8736, 32'd4287, -32'd1303},
{32'd3979, 32'd1133, -32'd5923, 32'd1390},
{32'd8767, 32'd12980, 32'd654, 32'd11195},
{-32'd816, -32'd18, 32'd2795, -32'd5172},
{-32'd2226, -32'd2521, 32'd7834, -32'd831},
{-32'd1665, 32'd327, -32'd4487, 32'd4342},
{-32'd6702, 32'd6130, -32'd4268, 32'd6831},
{-32'd8632, -32'd6505, 32'd5505, -32'd562},
{-32'd8572, -32'd4171, -32'd8583, 32'd3557},
{-32'd1686, -32'd2917, 32'd1067, -32'd7230},
{-32'd3976, 32'd7470, 32'd19303, 32'd2135},
{-32'd291, -32'd12743, 32'd3433, 32'd1435},
{-32'd14459, -32'd3277, 32'd2005, 32'd3158},
{-32'd128, 32'd8916, 32'd16529, -32'd7186},
{32'd14058, 32'd4809, 32'd19589, 32'd6466},
{32'd804, -32'd3429, 32'd790, -32'd2011},
{32'd382, -32'd8788, 32'd9382, -32'd3524},
{-32'd7556, -32'd7123, 32'd5536, -32'd6452},
{32'd4687, 32'd2589, -32'd5962, 32'd4672},
{32'd2111, -32'd4686, -32'd6274, -32'd11056},
{-32'd845, 32'd8338, 32'd5067, 32'd4449},
{-32'd2219, -32'd1602, -32'd4460, 32'd10998},
{32'd1443, 32'd6570, 32'd12493, 32'd368},
{-32'd5327, 32'd7936, -32'd5950, -32'd5894},
{32'd3714, 32'd7222, -32'd514, -32'd6058},
{-32'd2494, -32'd7263, -32'd4768, -32'd15748},
{-32'd8844, 32'd1284, -32'd11225, 32'd2039},
{32'd619, 32'd196, -32'd1722, 32'd6549},
{32'd6190, 32'd1567, -32'd15016, -32'd2879},
{32'd2699, -32'd11046, 32'd1733, -32'd12},
{32'd8268, 32'd1293, -32'd4229, -32'd5143},
{32'd13752, -32'd6441, 32'd8390, -32'd8366},
{-32'd19615, -32'd10472, 32'd11289, -32'd3287},
{-32'd5815, -32'd4485, -32'd14375, -32'd7819},
{-32'd9623, 32'd7590, 32'd9536, 32'd4429},
{32'd6150, -32'd6312, 32'd260, 32'd4979},
{-32'd803, 32'd5147, -32'd12930, 32'd10989},
{32'd96, 32'd12211, 32'd412, 32'd2958},
{32'd3646, 32'd1538, -32'd265, 32'd2520},
{-32'd5437, -32'd4199, 32'd13548, -32'd1214},
{-32'd3509, 32'd6342, -32'd2590, -32'd5995},
{-32'd15, -32'd4989, -32'd6979, 32'd6701},
{32'd6530, 32'd865, 32'd12698, -32'd6256},
{32'd5871, -32'd6205, -32'd10503, 32'd11577},
{-32'd1078, -32'd8775, -32'd3472, 32'd994},
{32'd1506, 32'd8167, -32'd5729, 32'd2670},
{32'd14537, -32'd2605, -32'd5177, 32'd3947},
{-32'd703, 32'd3959, -32'd518, -32'd5787},
{-32'd4047, -32'd13346, -32'd3784, -32'd3235},
{32'd1283, 32'd4963, -32'd16335, 32'd1491},
{32'd8211, 32'd1253, -32'd2306, -32'd9990},
{32'd3715, 32'd21217, 32'd14033, 32'd2985},
{-32'd3068, -32'd3736, 32'd2827, 32'd2500},
{-32'd4353, -32'd3758, 32'd2968, -32'd5602},
{-32'd4928, 32'd8468, -32'd10412, -32'd1326},
{32'd9350, -32'd11741, 32'd1608, 32'd5144},
{32'd28, -32'd446, -32'd5911, -32'd996},
{32'd8473, 32'd3317, 32'd5730, 32'd1146},
{-32'd8046, -32'd3884, 32'd1675, -32'd6416},
{32'd14216, -32'd7875, 32'd18731, -32'd84},
{32'd9235, 32'd8017, 32'd6389, 32'd7226},
{32'd5289, 32'd6767, -32'd4823, -32'd706},
{32'd20492, -32'd12567, -32'd5549, -32'd2163},
{32'd5385, -32'd10809, 32'd13884, 32'd6476},
{32'd3809, -32'd5112, 32'd880, -32'd2419},
{-32'd5089, 32'd2479, -32'd9965, 32'd2510},
{-32'd4878, 32'd2201, 32'd108, -32'd4009},
{32'd5734, -32'd1823, -32'd3605, -32'd7534},
{-32'd226, 32'd2677, -32'd1577, -32'd1955},
{-32'd958, -32'd1128, -32'd9685, -32'd5752},
{-32'd5225, -32'd5636, -32'd7810, 32'd9224},
{32'd4492, -32'd3812, -32'd6863, -32'd9487},
{-32'd2918, 32'd9455, 32'd1626, -32'd3762},
{-32'd1216, -32'd10369, -32'd283, 32'd1143},
{32'd5487, -32'd5811, -32'd6506, -32'd4071},
{32'd4332, -32'd7204, -32'd6284, -32'd1368},
{-32'd995, 32'd1523, 32'd9127, -32'd4544},
{32'd3015, -32'd10651, -32'd3608, 32'd2119},
{-32'd2916, -32'd2, 32'd1753, -32'd4299},
{32'd7284, 32'd4722, 32'd1415, -32'd8285},
{32'd3581, 32'd9319, 32'd7118, 32'd2067},
{-32'd9933, -32'd2612, 32'd25, 32'd1201},
{32'd1651, 32'd1379, -32'd12224, -32'd3161},
{-32'd897, 32'd4533, 32'd2984, 32'd8665},
{32'd268, -32'd611, 32'd10252, 32'd6750},
{32'd7341, 32'd7332, -32'd6156, 32'd11033},
{32'd6385, -32'd3003, 32'd3357, -32'd3287},
{32'd2073, -32'd4625, 32'd9193, -32'd15769},
{-32'd348, -32'd9524, 32'd2077, -32'd3684},
{32'd1742, 32'd219, -32'd3219, 32'd5254},
{32'd11540, -32'd1514, -32'd4056, 32'd2155},
{32'd7284, -32'd174, -32'd5317, -32'd1114},
{-32'd9956, -32'd3872, 32'd5345, -32'd8117},
{32'd8563, -32'd3122, 32'd1293, -32'd16223},
{32'd177, 32'd1059, 32'd37, 32'd4739},
{32'd10209, -32'd5184, -32'd8467, 32'd7780},
{32'd1963, -32'd7264, -32'd1370, 32'd2541},
{32'd2446, 32'd4219, -32'd2944, 32'd3001},
{32'd7334, 32'd289, 32'd2006, 32'd4004},
{32'd3246, 32'd4903, 32'd3188, 32'd2622},
{32'd2377, -32'd2119, -32'd7626, -32'd1126},
{32'd1901, 32'd1294, -32'd2919, 32'd4955},
{-32'd908, -32'd4169, 32'd2313, 32'd7112},
{-32'd6451, 32'd6808, 32'd1923, -32'd946},
{32'd12693, 32'd2051, 32'd1322, -32'd1264},
{32'd6838, 32'd3566, 32'd10846, 32'd3380},
{-32'd4091, 32'd1708, 32'd806, 32'd13497},
{32'd6563, -32'd2099, -32'd13974, -32'd919},
{-32'd2807, -32'd168, -32'd5408, 32'd6018},
{-32'd1869, 32'd4494, 32'd9596, 32'd369},
{-32'd11375, -32'd8244, -32'd1365, 32'd1911},
{32'd11286, -32'd1236, 32'd3266, 32'd2074},
{-32'd12975, -32'd3752, -32'd12009, 32'd6277},
{32'd9456, -32'd3372, -32'd1840, -32'd5383},
{32'd2507, -32'd5735, -32'd3328, -32'd10780},
{-32'd1068, -32'd2225, -32'd2249, 32'd7541},
{-32'd2361, 32'd6149, -32'd19697, 32'd4378},
{-32'd330, -32'd274, -32'd4539, -32'd2824},
{32'd2795, -32'd3823, 32'd1590, -32'd16935},
{-32'd5078, -32'd6607, 32'd9074, -32'd2468},
{32'd2754, 32'd7151, -32'd11482, -32'd4708},
{32'd3088, -32'd3899, -32'd12609, 32'd4140},
{32'd4867, 32'd8740, 32'd9, -32'd391},
{-32'd10476, 32'd2386, 32'd2875, 32'd5877},
{-32'd283, -32'd5035, 32'd10054, -32'd9843},
{-32'd3374, -32'd10419, -32'd2059, -32'd5125},
{-32'd8419, -32'd7720, 32'd3273, 32'd4438},
{-32'd7422, 32'd85, -32'd5388, 32'd1264},
{32'd11129, 32'd8448, 32'd7730, 32'd6313},
{32'd2304, 32'd82, 32'd7335, 32'd1979},
{32'd10197, 32'd8380, 32'd1343, 32'd2286},
{32'd9042, -32'd5952, 32'd9341, 32'd278},
{32'd3660, -32'd5968, -32'd10179, -32'd21042},
{-32'd468, -32'd18719, -32'd2312, 32'd2435},
{-32'd1894, 32'd8209, 32'd4049, -32'd1369},
{-32'd14346, -32'd11576, -32'd8579, -32'd6157},
{-32'd1681, -32'd1663, -32'd2148, -32'd5761},
{32'd4991, 32'd6164, -32'd920, 32'd7811},
{32'd3912, 32'd7233, -32'd833, -32'd2529},
{32'd6547, 32'd4265, -32'd7103, 32'd6170},
{-32'd10942, -32'd3452, 32'd6089, -32'd8043},
{-32'd747, 32'd629, -32'd4318, -32'd5345},
{-32'd7930, 32'd9434, 32'd5187, 32'd7165},
{-32'd5169, 32'd3133, 32'd1764, -32'd7646},
{32'd5635, 32'd1055, -32'd2505, -32'd17170},
{-32'd3830, 32'd4756, -32'd3911, -32'd7738},
{-32'd9566, -32'd3110, 32'd3884, -32'd7997},
{32'd2427, 32'd10855, -32'd693, 32'd12335},
{-32'd4335, 32'd8054, -32'd4943, 32'd1947},
{32'd26509, 32'd6549, -32'd2476, 32'd2510},
{-32'd1290, -32'd3189, 32'd14674, 32'd7694},
{-32'd5190, -32'd9488, 32'd5848, -32'd1538},
{-32'd455, -32'd2434, 32'd13111, -32'd3720},
{32'd7827, 32'd2857, -32'd9309, -32'd7544},
{32'd4711, 32'd5314, -32'd6306, -32'd9724},
{32'd1477, -32'd9947, -32'd14417, 32'd3684},
{-32'd14657, -32'd6871, 32'd7401, 32'd12041},
{-32'd14195, -32'd132, 32'd3839, -32'd11286},
{32'd328, 32'd7231, 32'd1337, 32'd3384},
{-32'd6301, 32'd6028, -32'd5382, -32'd8906},
{32'd249, -32'd4386, 32'd15864, -32'd45},
{32'd6536, -32'd3846, -32'd8380, -32'd5271},
{32'd110, 32'd8580, -32'd1209, -32'd12042},
{-32'd1290, 32'd6947, 32'd17482, 32'd3023},
{32'd5686, 32'd3896, 32'd5504, 32'd7654},
{32'd5979, -32'd10431, 32'd1350, -32'd8429},
{32'd6073, -32'd15629, -32'd1377, 32'd9077},
{32'd9845, -32'd4997, -32'd2293, -32'd12610},
{-32'd9195, -32'd3198, 32'd2013, 32'd13},
{32'd795, 32'd1174, -32'd10821, -32'd6811},
{-32'd6538, -32'd3857, -32'd1016, -32'd1715},
{-32'd5143, -32'd1597, -32'd19005, 32'd3059},
{-32'd1007, 32'd7712, 32'd9801, 32'd174},
{32'd9968, 32'd7494, -32'd2511, -32'd8304},
{32'd12855, 32'd2439, 32'd1588, -32'd756},
{32'd5163, -32'd9397, -32'd7305, 32'd5628},
{32'd3479, 32'd2419, -32'd1242, -32'd3081},
{32'd6205, -32'd12267, -32'd1933, -32'd1097},
{32'd9222, 32'd309, 32'd1012, -32'd2581},
{-32'd4860, 32'd8322, 32'd24770, -32'd784},
{32'd8886, 32'd7501, -32'd10596, -32'd2455},
{-32'd16068, -32'd5412, -32'd5224, -32'd1358},
{-32'd9129, 32'd1304, -32'd629, 32'd256},
{32'd11325, 32'd5709, 32'd2776, 32'd5684},
{-32'd1138, 32'd5063, 32'd1832, -32'd11050},
{-32'd7794, 32'd15374, -32'd6864, -32'd3150},
{-32'd4436, -32'd11945, -32'd2683, -32'd5385},
{32'd4432, -32'd2671, 32'd6432, -32'd3598},
{32'd2505, 32'd3004, 32'd5111, 32'd3993},
{32'd3192, 32'd91, 32'd5338, -32'd1300},
{32'd10079, -32'd4449, -32'd17567, -32'd9982},
{-32'd6697, -32'd10289, 32'd11719, 32'd1399},
{32'd15525, -32'd1662, -32'd732, 32'd6993},
{32'd1783, -32'd8469, -32'd5432, 32'd4379},
{-32'd1507, 32'd12821, 32'd2221, -32'd2696},
{32'd13568, 32'd13546, 32'd4228, 32'd5446},
{-32'd1054, -32'd4939, -32'd6645, -32'd7464},
{32'd3735, 32'd5104, -32'd14570, -32'd2382},
{-32'd7291, 32'd4292, -32'd6357, 32'd6934},
{-32'd3624, -32'd15082, -32'd1478, 32'd8377},
{-32'd844, -32'd3446, -32'd4303, -32'd10284},
{32'd6780, -32'd1291, -32'd11621, -32'd8769},
{-32'd4020, 32'd6513, -32'd4446, -32'd6356},
{-32'd2212, -32'd896, 32'd11781, -32'd1379},
{32'd6473, 32'd1133, -32'd1353, 32'd5262},
{-32'd7862, -32'd11603, -32'd7465, -32'd1692},
{32'd4834, 32'd3818, -32'd9599, -32'd5786},
{32'd11768, -32'd1162, 32'd6780, 32'd3575},
{32'd6642, 32'd8865, -32'd2138, -32'd2169},
{-32'd16361, -32'd2054, 32'd16432, -32'd714},
{32'd8447, -32'd4508, 32'd5243, -32'd1879},
{-32'd110, -32'd7558, 32'd7990, -32'd6035},
{32'd839, 32'd1088, -32'd494, -32'd8205},
{32'd11512, 32'd1519, -32'd13948, -32'd1518},
{-32'd7853, -32'd5207, -32'd1144, 32'd6613},
{32'd2492, 32'd4449, 32'd1392, -32'd205},
{-32'd10250, -32'd7986, -32'd3793, -32'd12368},
{32'd16168, 32'd13842, 32'd7894, -32'd8379},
{-32'd11026, -32'd734, 32'd3320, 32'd5343},
{32'd8443, 32'd2462, -32'd1096, 32'd10959},
{-32'd1459, -32'd6530, 32'd6453, -32'd18646},
{-32'd1849, -32'd3497, -32'd5368, -32'd4859},
{-32'd1872, -32'd3653, 32'd489, 32'd6811},
{-32'd546, -32'd7842, 32'd10742, -32'd2358},
{-32'd3897, 32'd1011, -32'd729, 32'd4060},
{32'd13490, -32'd5073, -32'd8839, -32'd1938},
{-32'd6857, 32'd927, 32'd5405, 32'd1968},
{32'd1628, 32'd7781, -32'd2874, 32'd5655},
{-32'd9305, -32'd9052, -32'd1974, 32'd2122},
{32'd8224, -32'd3768, 32'd11857, -32'd8378},
{32'd5832, 32'd11571, 32'd10333, 32'd6734},
{32'd850, -32'd3977, -32'd5750, -32'd871},
{-32'd6371, -32'd3198, -32'd5554, -32'd14316},
{-32'd5263, 32'd3451, -32'd6244, -32'd1080},
{-32'd2509, 32'd4228, 32'd20577, 32'd3071},
{32'd3546, -32'd1618, -32'd4086, 32'd4887},
{32'd7896, 32'd1104, 32'd4068, 32'd2677},
{32'd560, 32'd4673, 32'd3975, -32'd3201},
{32'd3597, -32'd296, 32'd824, -32'd3764},
{-32'd6745, -32'd12739, 32'd8487, -32'd644},
{32'd1115, -32'd3853, -32'd4451, -32'd2564},
{-32'd5058, 32'd5645, 32'd5281, -32'd1904},
{-32'd3731, 32'd1, -32'd3611, -32'd2926},
{32'd431, -32'd3266, -32'd3791, 32'd7676},
{-32'd5770, -32'd7076, 32'd5253, -32'd9124},
{-32'd6785, 32'd11528, 32'd4490, 32'd270},
{-32'd10644, 32'd7542, 32'd4086, -32'd3719},
{32'd10620, 32'd4708, -32'd6124, 32'd2950},
{-32'd1961, 32'd8146, -32'd11433, -32'd938},
{-32'd1304, 32'd1189, -32'd4961, 32'd1856},
{-32'd5703, 32'd8726, 32'd12197, -32'd119},
{-32'd7290, 32'd7187, 32'd2768, -32'd1865},
{32'd8980, 32'd3534, -32'd2293, -32'd2147},
{32'd5504, 32'd2884, -32'd182, 32'd2796},
{-32'd4723, -32'd9953, 32'd3468, 32'd6766},
{32'd9360, 32'd12445, 32'd3920, 32'd796},
{-32'd3773, 32'd4062, 32'd5633, 32'd1961},
{-32'd10862, 32'd12561, 32'd4123, -32'd13278},
{32'd6787, -32'd11443, 32'd6972, -32'd2404},
{-32'd627, 32'd3092, -32'd4736, 32'd2376},
{-32'd9354, 32'd4388, -32'd5554, -32'd4525},
{32'd320, -32'd9673, 32'd3747, 32'd9853},
{32'd6366, 32'd14485, 32'd7307, 32'd4507},
{-32'd5500, 32'd2181, 32'd6533, 32'd10422},
{-32'd7413, -32'd4744, -32'd4689, 32'd4674},
{-32'd8519, -32'd6119, 32'd582, -32'd4644},
{-32'd1650, 32'd5594, 32'd1432, -32'd2672},
{32'd11462, 32'd9391, -32'd12046, 32'd2714},
{32'd9460, 32'd3075, -32'd5915, 32'd6526},
{32'd5932, -32'd4980, -32'd711, -32'd6473},
{-32'd1713, 32'd5296, 32'd8645, 32'd8258},
{-32'd11447, -32'd5133, 32'd1030, -32'd15145},
{-32'd1579, 32'd6314, 32'd1720, 32'd13517},
{-32'd14571, -32'd2491, 32'd2616, -32'd6202},
{32'd5892, 32'd8558, -32'd5569, 32'd1713},
{32'd5427, -32'd8122, 32'd2320, 32'd8584},
{32'd4517, -32'd16188, 32'd4799, -32'd7524},
{32'd3837, 32'd4672, -32'd268, 32'd10172},
{-32'd14406, -32'd958, -32'd687, 32'd6074},
{-32'd4259, -32'd5402, 32'd4641, 32'd4065},
{32'd7093, -32'd4954, -32'd5551, -32'd4416},
{-32'd10102, -32'd5916, 32'd2828, -32'd2265},
{32'd2574, -32'd1243, -32'd1022, -32'd1203},
{-32'd4456, 32'd10502, -32'd687, 32'd6647},
{-32'd12553, -32'd2159, -32'd1691, 32'd4695},
{32'd4272, 32'd2305, -32'd15992, 32'd7816}
},
{{32'd4609, 32'd8492, 32'd1599, -32'd1288},
{-32'd2921, -32'd2369, -32'd3599, -32'd4628},
{32'd5333, 32'd1546, 32'd4307, 32'd6863},
{-32'd11689, 32'd2162, 32'd6990, -32'd10879},
{32'd9833, 32'd4779, -32'd4548, 32'd12524},
{-32'd1250, 32'd1632, 32'd7111, -32'd3731},
{-32'd6628, 32'd23, -32'd274, 32'd5185},
{-32'd440, -32'd6358, 32'd1745, -32'd8109},
{-32'd2888, -32'd3655, 32'd231, -32'd5564},
{32'd8952, 32'd11358, 32'd9417, 32'd1818},
{-32'd6739, -32'd5906, -32'd767, -32'd5238},
{32'd10059, -32'd11027, 32'd837, -32'd816},
{32'd7290, -32'd59, 32'd8375, -32'd1381},
{-32'd6642, -32'd94, 32'd872, -32'd833},
{-32'd13106, -32'd8484, -32'd4474, 32'd549},
{-32'd9147, -32'd1917, -32'd605, 32'd6558},
{-32'd3084, 32'd1196, -32'd218, -32'd4523},
{32'd9470, 32'd8577, -32'd1320, -32'd24},
{-32'd747, -32'd504, 32'd2481, 32'd6024},
{32'd4453, -32'd11965, 32'd4854, -32'd1388},
{32'd271, -32'd803, -32'd1453, 32'd1257},
{-32'd9266, 32'd1763, -32'd2968, 32'd2946},
{-32'd1206, -32'd1548, -32'd2625, 32'd1978},
{32'd1723, -32'd99, -32'd56, -32'd4941},
{32'd5700, 32'd1936, 32'd5735, 32'd3843},
{-32'd1812, 32'd2679, 32'd8149, -32'd3819},
{32'd2443, -32'd1839, -32'd7689, 32'd620},
{32'd5197, 32'd5984, -32'd248, -32'd1547},
{32'd3197, 32'd158, 32'd6944, 32'd13064},
{32'd2598, 32'd2723, 32'd3007, 32'd548},
{-32'd5699, -32'd2422, 32'd1978, 32'd3513},
{-32'd2357, -32'd6419, -32'd4874, -32'd5249},
{-32'd4772, -32'd26, -32'd306, 32'd3558},
{32'd1870, -32'd607, -32'd6105, 32'd3674},
{32'd11142, 32'd3418, 32'd5502, 32'd1671},
{-32'd2561, -32'd4198, 32'd4408, 32'd2128},
{32'd4730, 32'd1739, 32'd1906, -32'd3091},
{-32'd6857, -32'd973, -32'd3337, -32'd3435},
{-32'd3174, 32'd3548, 32'd490, 32'd658},
{32'd4792, 32'd1094, 32'd969, -32'd3784},
{32'd12840, 32'd6803, -32'd2106, -32'd3831},
{32'd3993, -32'd1091, 32'd5464, 32'd5641},
{32'd7012, 32'd3192, 32'd1746, -32'd650},
{-32'd6658, -32'd889, 32'd561, 32'd2796},
{-32'd706, 32'd1614, 32'd41, -32'd269},
{-32'd6850, 32'd7898, -32'd2732, -32'd1934},
{32'd2255, -32'd4642, 32'd685, -32'd4321},
{32'd1990, -32'd9101, -32'd4497, 32'd2009},
{-32'd3428, 32'd3031, 32'd3844, 32'd1490},
{-32'd1843, 32'd862, -32'd4816, -32'd2767},
{-32'd7092, -32'd8506, -32'd6311, -32'd3900},
{32'd7445, -32'd623, -32'd191, -32'd2915},
{-32'd1619, -32'd8656, -32'd3901, 32'd952},
{-32'd7370, -32'd1040, 32'd2653, 32'd391},
{32'd6454, 32'd3902, -32'd567, 32'd10346},
{-32'd5864, -32'd9682, -32'd3868, -32'd5110},
{32'd4684, -32'd5962, -32'd1812, 32'd8400},
{-32'd5788, -32'd3467, -32'd3073, 32'd3278},
{-32'd8416, 32'd446, -32'd2433, -32'd2805},
{32'd2278, -32'd4827, 32'd4378, 32'd10033},
{-32'd3669, -32'd2617, 32'd5264, 32'd1783},
{-32'd5093, -32'd3570, -32'd3251, 32'd1719},
{-32'd6447, -32'd10920, -32'd1717, -32'd7670},
{-32'd4645, -32'd4595, 32'd4307, 32'd8315},
{32'd7685, -32'd2192, -32'd684, -32'd2313},
{32'd9840, 32'd658, 32'd4683, 32'd3989},
{32'd10600, -32'd4781, 32'd1845, 32'd1814},
{32'd3628, -32'd7079, 32'd747, -32'd1926},
{32'd16873, 32'd2204, -32'd3712, -32'd7215},
{32'd5483, -32'd3207, 32'd102, -32'd9464},
{-32'd2597, -32'd6382, -32'd6878, 32'd498},
{32'd7561, 32'd7030, -32'd5284, 32'd3235},
{32'd4967, 32'd2691, -32'd1982, 32'd6686},
{32'd3386, -32'd1521, -32'd3795, -32'd4983},
{32'd3390, 32'd11682, 32'd2859, 32'd7886},
{32'd8804, 32'd1892, 32'd5577, -32'd8242},
{-32'd899, -32'd1525, -32'd6085, -32'd12421},
{32'd1910, 32'd1528, -32'd3685, 32'd2575},
{32'd1586, 32'd3777, 32'd6064, -32'd3881},
{-32'd6287, 32'd2853, 32'd2063, 32'd435},
{-32'd3820, 32'd1604, 32'd3427, -32'd2683},
{32'd2926, -32'd212, 32'd8500, 32'd626},
{32'd218, 32'd1853, -32'd4919, -32'd4069},
{-32'd5406, -32'd4477, -32'd8383, 32'd2657},
{32'd7594, -32'd7346, -32'd4707, -32'd3103},
{-32'd7902, -32'd4612, -32'd7468, 32'd7906},
{-32'd180, -32'd335, 32'd2295, 32'd3836},
{-32'd734, -32'd1604, -32'd8446, -32'd2960},
{32'd4262, -32'd5543, -32'd2342, 32'd2711},
{-32'd7937, -32'd1090, -32'd2893, -32'd420},
{-32'd523, 32'd5859, 32'd6158, -32'd4622},
{-32'd6346, -32'd3265, -32'd4397, -32'd411},
{32'd3322, 32'd7485, 32'd5641, 32'd3919},
{32'd5462, -32'd1582, 32'd6953, 32'd2454},
{-32'd3863, 32'd3441, 32'd1234, 32'd823},
{-32'd2387, -32'd2087, 32'd655, -32'd11621},
{-32'd6332, 32'd8971, 32'd8184, -32'd1536},
{32'd3834, 32'd3033, 32'd2162, -32'd1693},
{32'd133, 32'd330, -32'd683, 32'd4785},
{32'd6091, 32'd12599, 32'd7897, 32'd4408},
{-32'd1339, 32'd4071, 32'd7468, -32'd5827},
{32'd1986, -32'd714, -32'd553, -32'd4621},
{32'd286, -32'd4499, 32'd3007, -32'd12690},
{32'd2799, -32'd2359, -32'd5541, -32'd8825},
{32'd4201, 32'd7271, -32'd4715, 32'd546},
{-32'd16949, 32'd6920, 32'd2761, 32'd5462},
{32'd6204, -32'd2585, 32'd5934, -32'd970},
{-32'd16821, -32'd1361, -32'd8191, 32'd2863},
{32'd7039, 32'd4577, 32'd6198, 32'd3678},
{32'd9507, -32'd4310, -32'd1168, 32'd5687},
{32'd9985, -32'd3901, -32'd7033, -32'd3005},
{32'd5524, 32'd2558, 32'd404, -32'd2134},
{32'd1515, 32'd4297, 32'd4548, 32'd104},
{32'd8881, 32'd2806, -32'd1137, -32'd4074},
{-32'd7902, 32'd1486, 32'd9163, -32'd258},
{32'd6200, -32'd892, -32'd385, 32'd4798},
{-32'd3799, 32'd3936, 32'd6620, 32'd8187},
{32'd1871, -32'd3097, -32'd2228, -32'd9561},
{-32'd4989, -32'd7600, -32'd3945, 32'd3067},
{-32'd196, 32'd6583, 32'd9482, 32'd3620},
{-32'd1783, 32'd7458, 32'd9999, 32'd2111},
{32'd339, 32'd9814, -32'd6114, 32'd2052},
{32'd4352, 32'd2850, -32'd1683, 32'd6288},
{-32'd1627, -32'd253, 32'd4629, -32'd6438},
{-32'd5341, 32'd1641, -32'd1278, -32'd1802},
{32'd5815, 32'd5609, 32'd5347, -32'd10387},
{-32'd3500, 32'd5435, 32'd2370, -32'd4856},
{-32'd1579, -32'd1421, -32'd780, -32'd4392},
{-32'd4472, -32'd1832, 32'd2437, -32'd1613},
{32'd1008, 32'd188, -32'd10535, 32'd2548},
{32'd10317, -32'd2185, -32'd4369, 32'd4267},
{32'd3072, -32'd1803, -32'd931, -32'd8126},
{-32'd8112, -32'd2413, -32'd2569, 32'd1472},
{32'd5040, 32'd1756, 32'd2659, 32'd4702},
{-32'd6356, 32'd2095, 32'd141, 32'd1572},
{-32'd10127, -32'd5263, -32'd8631, -32'd914},
{32'd155, 32'd1033, 32'd6360, 32'd1069},
{-32'd1443, 32'd1202, 32'd3661, -32'd6077},
{32'd7720, 32'd3630, 32'd3458, -32'd2347},
{32'd973, 32'd228, -32'd6061, -32'd7928},
{-32'd7, -32'd3965, -32'd3473, -32'd7364},
{-32'd9146, -32'd8562, 32'd3761, -32'd4688},
{-32'd5964, -32'd2689, -32'd1805, 32'd2641},
{-32'd5036, 32'd264, -32'd266, -32'd3437},
{32'd8960, 32'd4159, 32'd5778, 32'd2898},
{32'd13784, -32'd6774, 32'd3105, -32'd3702},
{32'd728, 32'd3958, -32'd3442, 32'd1455},
{32'd1535, 32'd1526, 32'd409, 32'd2114},
{32'd2542, 32'd758, -32'd1746, 32'd3430},
{32'd5815, -32'd1546, -32'd439, -32'd2910},
{-32'd6954, -32'd828, -32'd5428, 32'd623},
{32'd1635, 32'd10134, -32'd3865, 32'd5271},
{-32'd11321, 32'd3610, -32'd3208, 32'd6837},
{32'd5665, 32'd5121, 32'd3329, 32'd1752},
{-32'd4767, -32'd13160, -32'd2652, -32'd6653},
{-32'd10675, 32'd10760, -32'd1570, 32'd6954},
{32'd5673, 32'd8341, 32'd2911, 32'd4808},
{-32'd1088, 32'd2314, -32'd3548, 32'd554},
{-32'd13172, 32'd4176, -32'd7337, 32'd6224},
{32'd10679, 32'd5886, 32'd5800, 32'd671},
{32'd3812, -32'd3677, -32'd653, -32'd3338},
{32'd11002, 32'd9773, 32'd10928, 32'd5795},
{32'd8323, -32'd4137, -32'd4408, -32'd3956},
{32'd1706, 32'd7728, -32'd583, -32'd4519},
{32'd5672, 32'd4160, 32'd1071, 32'd3712},
{-32'd4428, -32'd3664, -32'd3984, -32'd11432},
{32'd1085, -32'd2212, 32'd1803, 32'd5892},
{-32'd1257, -32'd5981, -32'd4696, -32'd176},
{-32'd7322, -32'd71, -32'd4120, 32'd2953},
{-32'd12322, -32'd5875, -32'd6233, 32'd3825},
{32'd2640, -32'd3255, -32'd7513, -32'd1639},
{32'd3152, -32'd4219, -32'd2046, -32'd4419},
{32'd7552, 32'd3097, 32'd5413, -32'd2754},
{-32'd1378, -32'd4006, -32'd2684, -32'd3665},
{-32'd12125, -32'd1836, -32'd5386, -32'd4140},
{32'd1027, 32'd3986, -32'd2912, 32'd5771},
{-32'd2927, 32'd2466, 32'd160, -32'd3110},
{-32'd5369, 32'd1152, -32'd5062, -32'd6518},
{-32'd3621, 32'd954, 32'd1494, 32'd5003},
{-32'd4821, -32'd5094, 32'd713, 32'd773},
{32'd108, -32'd7552, -32'd2253, -32'd2190},
{-32'd10066, 32'd3473, -32'd3205, 32'd626},
{-32'd3313, -32'd5008, -32'd783, -32'd2439},
{32'd3833, 32'd6901, -32'd3588, 32'd2324},
{-32'd3894, -32'd3168, 32'd8043, -32'd2364},
{-32'd3739, -32'd2308, 32'd128, -32'd1199},
{32'd2494, -32'd3944, 32'd11459, 32'd4407},
{-32'd1129, 32'd8587, -32'd3035, -32'd2608},
{-32'd10776, -32'd1206, 32'd2376, -32'd2175},
{-32'd11261, 32'd2158, -32'd4397, 32'd5253},
{-32'd2697, 32'd2235, 32'd3408, 32'd2830},
{-32'd4848, -32'd12729, -32'd4974, -32'd5272},
{-32'd3962, -32'd3043, 32'd1552, -32'd1598},
{32'd2831, 32'd6513, -32'd716, 32'd7255},
{32'd5202, -32'd732, -32'd1546, -32'd1934},
{-32'd796, 32'd5485, 32'd3957, 32'd4658},
{32'd7711, 32'd1671, -32'd8447, 32'd832},
{-32'd1175, -32'd43, -32'd10319, 32'd682},
{32'd4251, 32'd345, -32'd4479, 32'd2352},
{32'd4532, -32'd445, 32'd6271, -32'd5574},
{-32'd3329, -32'd8565, -32'd6636, -32'd4314},
{32'd10343, 32'd2786, -32'd174, -32'd3730},
{32'd4716, -32'd847, -32'd3070, -32'd4633},
{32'd7568, -32'd9596, -32'd5506, -32'd1653},
{32'd3699, -32'd11319, -32'd2453, -32'd5812},
{32'd6588, 32'd1385, -32'd354, -32'd6847},
{32'd2928, 32'd14047, 32'd2727, 32'd1972},
{-32'd6005, -32'd6202, -32'd5236, -32'd8846},
{-32'd6297, 32'd1450, 32'd6824, 32'd5173},
{32'd1711, 32'd8978, -32'd2412, 32'd4618},
{32'd3674, -32'd2400, 32'd3708, 32'd6977},
{-32'd401, -32'd305, 32'd1005, 32'd5337},
{-32'd612, -32'd4044, -32'd2116, -32'd4120},
{32'd5048, 32'd7787, -32'd472, -32'd5930},
{32'd10492, 32'd4484, 32'd1012, 32'd976},
{-32'd12537, 32'd2551, -32'd2871, -32'd1075},
{32'd3757, -32'd7487, 32'd6422, -32'd9936},
{-32'd3784, 32'd257, -32'd4006, 32'd1211},
{-32'd5718, -32'd1613, 32'd2607, 32'd2495},
{32'd30, 32'd7565, -32'd341, -32'd4545},
{-32'd1347, -32'd3997, 32'd2323, -32'd7497},
{32'd745, 32'd6655, 32'd3304, 32'd6128},
{-32'd11200, 32'd5776, 32'd7498, 32'd2198},
{32'd2114, 32'd2268, 32'd805, 32'd3812},
{-32'd1008, -32'd1068, 32'd996, 32'd18450},
{-32'd4520, -32'd1695, 32'd1002, -32'd2155},
{32'd1840, -32'd8293, -32'd906, -32'd4989},
{-32'd862, -32'd1397, 32'd4754, 32'd2781},
{32'd10760, -32'd9934, 32'd51, -32'd2251},
{32'd7538, 32'd2039, 32'd4145, -32'd3620},
{-32'd4044, -32'd2687, -32'd5174, 32'd6276},
{32'd7382, -32'd2825, -32'd2716, -32'd9126},
{-32'd2361, 32'd3653, 32'd1268, 32'd2758},
{32'd7871, 32'd5307, 32'd947, 32'd1572},
{-32'd4054, -32'd5076, -32'd1283, -32'd8439},
{32'd5068, -32'd403, 32'd5965, -32'd7562},
{32'd187, -32'd113, -32'd3811, 32'd6095},
{-32'd4345, 32'd6816, -32'd1074, -32'd1869},
{-32'd4698, 32'd3553, -32'd4315, 32'd6343},
{32'd1269, 32'd2285, -32'd2354, 32'd5564},
{32'd7019, 32'd6853, 32'd711, 32'd3331},
{-32'd4015, 32'd1736, -32'd7187, -32'd1510},
{-32'd15100, -32'd6516, -32'd6333, -32'd236},
{-32'd2678, -32'd6520, -32'd3672, -32'd988},
{-32'd864, 32'd9439, 32'd7658, 32'd1144},
{32'd2939, -32'd2931, -32'd1389, -32'd889},
{32'd5830, -32'd1136, -32'd4147, 32'd6504},
{32'd11792, -32'd1685, 32'd1931, -32'd921},
{-32'd3577, 32'd6707, 32'd3503, -32'd3014},
{-32'd15798, 32'd220, 32'd3712, -32'd590},
{-32'd230, -32'd6615, 32'd2937, 32'd14588},
{32'd3452, -32'd116, 32'd3781, -32'd4863},
{32'd10247, 32'd3719, 32'd5156, 32'd8132},
{-32'd4846, -32'd8715, 32'd1691, -32'd5227},
{-32'd11345, 32'd950, -32'd9453, -32'd8723},
{-32'd1182, -32'd5062, 32'd2046, -32'd3183},
{32'd938, -32'd8178, 32'd4615, -32'd2686},
{32'd9146, 32'd2522, 32'd1787, -32'd7466},
{-32'd4038, -32'd870, -32'd10395, -32'd1590},
{32'd7516, 32'd4443, 32'd4058, -32'd4477},
{-32'd2848, -32'd3823, 32'd3412, -32'd3897},
{32'd9651, -32'd495, 32'd815, 32'd8187},
{-32'd3811, 32'd2696, 32'd1567, -32'd2734},
{32'd1337, 32'd1559, -32'd3428, -32'd8923},
{32'd5945, 32'd1873, -32'd1138, -32'd618},
{-32'd2663, -32'd1759, 32'd867, -32'd6509},
{-32'd2863, 32'd5221, 32'd4152, -32'd4283},
{32'd1704, 32'd2182, -32'd7478, 32'd7805},
{-32'd4767, -32'd4972, -32'd7611, -32'd7557},
{32'd1799, -32'd7815, -32'd1028, 32'd4449},
{32'd4943, -32'd2014, -32'd2199, -32'd60},
{32'd7970, 32'd2861, -32'd816, 32'd10295},
{-32'd9985, -32'd3879, 32'd625, -32'd5819},
{32'd1398, -32'd2518, 32'd1663, 32'd4974},
{-32'd2108, -32'd1993, -32'd1158, 32'd3970},
{-32'd1700, -32'd8953, -32'd398, 32'd2915},
{32'd10134, 32'd13120, 32'd6656, 32'd3312},
{32'd6911, -32'd4128, 32'd1778, 32'd1432},
{-32'd7146, -32'd7558, -32'd7548, 32'd4844},
{-32'd6668, 32'd1082, -32'd8245, -32'd784},
{-32'd1514, 32'd4158, 32'd2725, 32'd4357},
{32'd8743, 32'd1631, 32'd1977, -32'd5177},
{32'd5107, 32'd3480, 32'd3115, 32'd2025},
{-32'd6556, -32'd3934, -32'd2928, -32'd3911},
{32'd364, 32'd1807, 32'd2799, 32'd2009},
{-32'd1751, -32'd7734, -32'd6988, 32'd164},
{32'd9200, 32'd5809, -32'd56, -32'd21},
{32'd3651, 32'd5378, -32'd5873, 32'd1331},
{-32'd1720, -32'd905, 32'd592, 32'd17529},
{-32'd4085, -32'd1649, -32'd8023, 32'd3221},
{-32'd5999, 32'd5021, 32'd8223, 32'd3511},
{-32'd4439, 32'd11575, 32'd4901, 32'd3939},
{32'd7533, 32'd8597, -32'd5862, 32'd2799},
{32'd6870, 32'd2866, -32'd7098, -32'd9187},
{-32'd8672, 32'd1953, -32'd8825, -32'd4490},
{-32'd8201, -32'd7286, -32'd1662, 32'd3344},
{32'd1907, -32'd2971, 32'd4146, -32'd2234},
{32'd741, 32'd6197, 32'd2638, -32'd842},
{32'd5492, 32'd620, 32'd5686, -32'd2674},
{32'd1501, 32'd1643, -32'd7072, -32'd1170}
},
{{-32'd192, 32'd6347, 32'd1860, 32'd3411},
{-32'd2421, 32'd7261, -32'd9405, -32'd5749},
{-32'd4754, 32'd6301, -32'd8974, 32'd1379},
{32'd1357, 32'd5827, 32'd1893, 32'd7039},
{32'd8790, 32'd1656, -32'd4663, -32'd394},
{-32'd8238, -32'd1860, -32'd9333, 32'd3684},
{-32'd2906, 32'd6796, 32'd5692, -32'd2888},
{-32'd8991, 32'd4783, -32'd156, 32'd6580},
{32'd4319, -32'd434, -32'd4612, -32'd2265},
{32'd8494, 32'd6182, -32'd1404, 32'd11852},
{-32'd2207, -32'd13356, -32'd1080, 32'd1624},
{-32'd7786, -32'd8124, -32'd16546, 32'd8795},
{32'd67, 32'd1992, 32'd3240, -32'd2410},
{-32'd16734, -32'd5751, -32'd3248, -32'd971},
{-32'd6090, -32'd9155, 32'd5577, 32'd84},
{-32'd3730, 32'd5404, 32'd7418, -32'd9386},
{32'd7136, 32'd3226, 32'd3765, 32'd8786},
{32'd732, -32'd8754, 32'd17982, -32'd4550},
{-32'd2752, -32'd7857, -32'd1418, 32'd3436},
{-32'd367, -32'd7739, -32'd5458, -32'd619},
{32'd3598, 32'd5615, -32'd3584, -32'd1773},
{-32'd2963, 32'd2407, 32'd1526, -32'd2214},
{-32'd1871, 32'd3065, -32'd5496, -32'd4832},
{-32'd13043, -32'd8279, 32'd7642, -32'd4311},
{-32'd1299, 32'd272, -32'd1867, 32'd13120},
{-32'd6025, 32'd2230, 32'd2105, -32'd9273},
{-32'd757, -32'd14270, -32'd5639, -32'd390},
{-32'd2862, 32'd8370, 32'd1592, -32'd602},
{32'd5109, 32'd6167, 32'd3445, 32'd516},
{-32'd2151, -32'd6923, 32'd11809, -32'd4066},
{-32'd17664, -32'd849, -32'd5861, 32'd8399},
{-32'd10927, -32'd1165, 32'd3822, -32'd270},
{32'd5157, 32'd2823, -32'd370, 32'd6003},
{-32'd10458, 32'd869, 32'd4902, -32'd8522},
{32'd3894, 32'd3837, 32'd373, 32'd964},
{-32'd1173, -32'd6515, -32'd6896, -32'd417},
{-32'd4309, -32'd2837, -32'd8004, 32'd14051},
{-32'd2717, -32'd6629, -32'd5960, -32'd222},
{32'd13211, -32'd10324, 32'd5934, -32'd4312},
{-32'd1456, -32'd5584, 32'd12507, 32'd1524},
{-32'd4253, -32'd253, -32'd6608, -32'd130},
{32'd6621, 32'd3213, 32'd7658, -32'd3145},
{32'd8094, 32'd3329, -32'd2699, 32'd6602},
{-32'd9068, -32'd484, -32'd242, -32'd9066},
{-32'd1997, -32'd5973, -32'd628, -32'd6103},
{32'd7969, -32'd11527, 32'd4234, -32'd3504},
{-32'd2672, -32'd7073, -32'd2656, -32'd5618},
{-32'd14142, -32'd2743, 32'd11484, -32'd3643},
{32'd7727, 32'd524, 32'd3368, 32'd3801},
{32'd1843, 32'd1747, -32'd4420, 32'd2170},
{-32'd2222, 32'd677, -32'd2896, -32'd3509},
{-32'd323, -32'd5628, -32'd882, 32'd951},
{-32'd2052, -32'd1108, -32'd6649, -32'd5632},
{32'd6880, 32'd1240, -32'd6, 32'd2985},
{-32'd5718, -32'd1223, 32'd4799, -32'd645},
{32'd153, -32'd1670, 32'd2907, 32'd3866},
{32'd479, -32'd2143, 32'd14773, -32'd2938},
{-32'd15768, 32'd7827, 32'd6906, -32'd5296},
{-32'd9231, -32'd3471, 32'd8053, 32'd7766},
{-32'd1007, 32'd2210, 32'd1903, -32'd3712},
{-32'd1227, -32'd15712, -32'd9665, 32'd2244},
{32'd901, 32'd2576, 32'd7327, -32'd3270},
{-32'd15343, -32'd6510, 32'd1784, -32'd3629},
{32'd3034, 32'd4083, -32'd3935, 32'd7296},
{32'd7598, 32'd2657, -32'd4516, -32'd5156},
{32'd2977, 32'd1771, 32'd10621, 32'd3369},
{32'd4936, -32'd9430, -32'd14124, 32'd14523},
{-32'd6723, -32'd11036, -32'd7358, -32'd7220},
{-32'd372, -32'd3314, 32'd7069, -32'd4455},
{-32'd557, 32'd4120, 32'd8341, -32'd4534},
{-32'd264, -32'd2216, 32'd6678, 32'd8455},
{-32'd2359, 32'd7776, 32'd6152, -32'd7701},
{-32'd10857, -32'd7298, 32'd6881, -32'd5340},
{32'd4815, -32'd7774, 32'd4620, 32'd1442},
{32'd6195, 32'd7119, 32'd4699, 32'd3103},
{-32'd2272, -32'd967, -32'd5008, -32'd9642},
{-32'd3687, 32'd698, 32'd3336, -32'd7080},
{-32'd5011, -32'd11348, -32'd1405, -32'd6553},
{32'd3636, 32'd2738, 32'd7131, -32'd1990},
{32'd6959, 32'd9457, 32'd10486, 32'd799},
{32'd5145, -32'd309, -32'd7991, 32'd7430},
{32'd3802, 32'd2572, -32'd916, 32'd1176},
{-32'd6014, 32'd8606, -32'd1643, 32'd1768},
{-32'd2871, 32'd10194, -32'd575, 32'd8377},
{32'd3133, 32'd2554, 32'd7141, -32'd11165},
{-32'd1739, -32'd4574, -32'd9237, -32'd2449},
{-32'd2711, 32'd2607, 32'd96, -32'd2041},
{-32'd7503, -32'd12718, 32'd22, -32'd2480},
{32'd1312, 32'd6053, 32'd287, -32'd3797},
{-32'd7389, -32'd4833, -32'd8023, 32'd4552},
{32'd1605, 32'd10754, 32'd2421, 32'd1543},
{-32'd4308, -32'd16679, -32'd4710, -32'd7072},
{-32'd2510, 32'd62, -32'd4928, -32'd2128},
{32'd4826, 32'd6373, -32'd6716, 32'd9478},
{32'd5317, 32'd1003, 32'd6925, 32'd1728},
{-32'd3314, 32'd490, -32'd10278, 32'd479},
{32'd10948, 32'd5984, 32'd2835, -32'd9106},
{-32'd1230, 32'd8765, 32'd5047, 32'd737},
{32'd506, -32'd424, -32'd1201, -32'd10084},
{32'd8121, 32'd9617, 32'd7530, -32'd1678},
{32'd1268, 32'd3255, -32'd13634, -32'd3375},
{-32'd9925, -32'd5486, 32'd5947, -32'd4933},
{32'd3686, 32'd5976, 32'd8070, 32'd3353},
{32'd3022, 32'd3315, 32'd1744, -32'd483},
{-32'd12084, 32'd6490, 32'd8081, -32'd190},
{32'd7028, 32'd6429, -32'd12409, 32'd2070},
{-32'd6431, -32'd1, -32'd7061, 32'd4855},
{-32'd5117, 32'd6434, -32'd5056, 32'd5610},
{-32'd6890, -32'd11379, 32'd719, -32'd2622},
{-32'd5317, -32'd4982, 32'd681, -32'd9491},
{32'd3887, -32'd5286, -32'd4820, -32'd4586},
{32'd11351, 32'd481, 32'd4697, 32'd2333},
{32'd4213, 32'd6585, -32'd155, 32'd14172},
{32'd8438, -32'd6960, -32'd11354, -32'd10033},
{-32'd4789, -32'd3515, -32'd6938, -32'd3468},
{32'd8635, 32'd260, -32'd5670, 32'd11363},
{-32'd2077, 32'd5954, -32'd5077, -32'd3825},
{32'd4194, -32'd12302, 32'd1108, 32'd3812},
{-32'd5247, 32'd5414, 32'd2844, 32'd7278},
{32'd800, 32'd7203, -32'd6901, 32'd7282},
{-32'd13408, -32'd12426, -32'd11097, 32'd3744},
{32'd5778, -32'd3592, -32'd8494, 32'd537},
{32'd8499, -32'd749, -32'd8316, -32'd449},
{-32'd5225, 32'd410, -32'd1368, 32'd5769},
{32'd4706, 32'd8494, -32'd4283, -32'd3954},
{32'd1332, -32'd7924, -32'd3898, -32'd6173},
{-32'd3073, 32'd905, -32'd171, -32'd2931},
{-32'd6138, -32'd8112, 32'd3744, -32'd2481},
{32'd3874, 32'd444, -32'd2011, -32'd2248},
{-32'd663, 32'd3218, 32'd4490, -32'd11624},
{32'd2825, 32'd2946, -32'd2773, -32'd4814},
{-32'd3528, 32'd687, -32'd751, -32'd8673},
{-32'd13458, -32'd11994, 32'd3441, 32'd604},
{32'd1202, 32'd5002, -32'd2642, 32'd4044},
{-32'd7925, -32'd7210, -32'd572, 32'd7258},
{32'd8022, 32'd3589, 32'd7428, 32'd10084},
{32'd10495, -32'd1631, 32'd1872, -32'd2512},
{32'd2921, -32'd7096, -32'd16425, -32'd4361},
{32'd1858, 32'd19726, -32'd6819, 32'd3822},
{32'd215, -32'd1991, -32'd6699, -32'd195},
{32'd2891, -32'd4064, -32'd273, 32'd665},
{-32'd9501, -32'd952, 32'd5023, -32'd2864},
{32'd5284, 32'd4550, 32'd14946, 32'd6082},
{-32'd11455, 32'd10676, -32'd6049, 32'd2682},
{32'd4994, -32'd4429, -32'd7822, 32'd6061},
{32'd13083, -32'd2094, -32'd3046, 32'd2130},
{-32'd5976, 32'd1383, -32'd5017, -32'd625},
{-32'd6121, -32'd12030, -32'd2775, 32'd2042},
{32'd3038, 32'd3539, 32'd2429, -32'd2816},
{-32'd18226, -32'd6392, -32'd10161, -32'd9136},
{-32'd6752, -32'd4541, 32'd934, -32'd4034},
{32'd4597, 32'd7829, -32'd7219, 32'd15059},
{32'd482, 32'd7579, -32'd4209, -32'd2556},
{-32'd6458, -32'd2970, 32'd1266, -32'd3615},
{-32'd14223, -32'd19691, 32'd3429, -32'd2870},
{32'd3032, 32'd13409, 32'd3564, -32'd3795},
{32'd3871, 32'd5829, -32'd8815, 32'd2935},
{32'd3304, -32'd9767, -32'd1300, 32'd5195},
{-32'd4611, 32'd355, -32'd2704, 32'd966},
{32'd2506, -32'd548, -32'd1965, -32'd868},
{-32'd3279, 32'd2455, 32'd8724, -32'd398},
{32'd3384, 32'd656, -32'd14357, -32'd1072},
{-32'd4069, -32'd16769, -32'd4157, 32'd2855},
{32'd5000, 32'd17299, 32'd5733, 32'd11582},
{32'd3432, 32'd11712, 32'd8460, -32'd8562},
{-32'd6495, -32'd6787, 32'd6228, 32'd5607},
{-32'd3052, 32'd4854, -32'd794, 32'd893},
{-32'd2015, -32'd3908, 32'd3443, -32'd3122},
{32'd778, -32'd5325, 32'd12607, -32'd8684},
{-32'd3145, 32'd5567, -32'd1822, -32'd14986},
{-32'd7786, -32'd7550, 32'd8781, -32'd1047},
{-32'd7647, -32'd970, -32'd1900, 32'd8859},
{32'd4088, 32'd7941, 32'd6452, 32'd7822},
{-32'd4478, -32'd9840, -32'd5500, 32'd2342},
{32'd1027, 32'd799, 32'd8707, -32'd6333},
{-32'd3902, 32'd10268, 32'd3367, -32'd6723},
{32'd9568, -32'd1946, 32'd7298, 32'd11279},
{-32'd3701, -32'd5791, -32'd8820, 32'd6968},
{-32'd4633, 32'd14643, 32'd8226, 32'd2720},
{-32'd1849, 32'd1183, -32'd1557, -32'd2739},
{-32'd6594, -32'd6233, 32'd2019, 32'd8096},
{-32'd6160, 32'd2254, 32'd453, -32'd1153},
{-32'd5872, -32'd8187, 32'd593, -32'd3176},
{-32'd3733, -32'd6050, 32'd1884, 32'd10490},
{-32'd10902, 32'd4249, -32'd4111, 32'd3369},
{32'd7751, 32'd3745, -32'd1654, 32'd3565},
{32'd6479, 32'd13477, 32'd2798, -32'd8149},
{-32'd2158, 32'd6639, -32'd1321, 32'd7033},
{32'd670, -32'd1423, 32'd8708, 32'd9707},
{32'd4354, 32'd6109, 32'd4378, 32'd1048},
{-32'd170, -32'd1359, -32'd12760, 32'd3197},
{-32'd8164, -32'd1787, 32'd6784, -32'd14226},
{-32'd6416, -32'd4982, 32'd3862, 32'd958},
{-32'd12592, -32'd1886, 32'd264, 32'd2817},
{-32'd11434, 32'd2540, -32'd8462, -32'd3533},
{-32'd5815, -32'd11419, -32'd11548, -32'd3815},
{-32'd3458, -32'd16012, -32'd7847, 32'd3316},
{32'd5529, -32'd7074, -32'd3212, 32'd5307},
{-32'd3807, -32'd2934, 32'd3445, 32'd6556},
{32'd11932, -32'd2973, -32'd2778, 32'd7867},
{-32'd5433, -32'd8353, 32'd1989, -32'd2051},
{-32'd6345, -32'd10130, -32'd11870, 32'd6157},
{32'd2498, 32'd13154, 32'd630, 32'd6766},
{32'd2508, 32'd5699, 32'd3093, 32'd9747},
{-32'd2351, 32'd11437, -32'd10511, 32'd6125},
{-32'd1996, -32'd790, 32'd3478, 32'd2542},
{-32'd4027, 32'd9332, 32'd780, 32'd2427},
{-32'd1917, -32'd5215, 32'd6855, 32'd1017},
{-32'd12993, 32'd4998, 32'd4669, -32'd10204},
{32'd1064, 32'd97, 32'd2967, -32'd3919},
{-32'd3254, -32'd7341, -32'd6250, -32'd2212},
{-32'd9242, -32'd10361, -32'd11796, 32'd3579},
{32'd3028, -32'd7308, -32'd6833, -32'd1387},
{-32'd1696, -32'd8595, 32'd5845, -32'd1850},
{-32'd516, -32'd14992, -32'd4598, 32'd650},
{-32'd3782, 32'd6814, -32'd784, 32'd2730},
{-32'd3397, -32'd4464, 32'd3692, 32'd13886},
{-32'd10488, 32'd1839, 32'd3772, -32'd390},
{32'd7209, 32'd10181, 32'd6711, 32'd7082},
{32'd1143, 32'd15089, 32'd10432, -32'd5936},
{-32'd9479, 32'd2809, 32'd7196, -32'd2436},
{-32'd543, -32'd77, -32'd5258, -32'd7901},
{32'd3163, -32'd615, -32'd2735, 32'd6780},
{-32'd4788, -32'd3333, 32'd13173, -32'd6736},
{-32'd5101, -32'd1289, -32'd8863, -32'd16234},
{32'd9579, 32'd15973, 32'd3746, -32'd2725},
{32'd6497, 32'd7014, 32'd2488, 32'd8026},
{32'd5761, 32'd2554, 32'd934, 32'd761},
{32'd4077, 32'd8162, -32'd5183, -32'd7039},
{32'd2320, -32'd5128, -32'd1297, 32'd8673},
{32'd541, -32'd3393, 32'd7, -32'd10894},
{32'd5, -32'd17757, 32'd2185, -32'd4058},
{-32'd1540, -32'd3326, -32'd6998, 32'd284},
{32'd2159, 32'd3748, -32'd7184, -32'd11963},
{32'd4051, 32'd2080, -32'd1226, -32'd1110},
{-32'd10493, -32'd13893, -32'd8281, -32'd3064},
{-32'd11474, 32'd14225, 32'd5651, -32'd7654},
{-32'd1198, -32'd13500, -32'd3472, 32'd3385},
{-32'd3362, -32'd5847, 32'd12945, -32'd2928},
{32'd2018, 32'd9925, 32'd4838, -32'd2962},
{32'd2288, -32'd8196, -32'd1439, 32'd1095},
{32'd202, 32'd3707, -32'd2643, -32'd3797},
{-32'd16940, -32'd12842, -32'd4495, -32'd7308},
{-32'd7413, -32'd8016, 32'd969, 32'd6733},
{32'd11707, 32'd3435, -32'd5389, 32'd2623},
{32'd4161, 32'd1114, 32'd7615, -32'd3965},
{-32'd9842, 32'd6110, 32'd2677, -32'd4066},
{-32'd1100, -32'd10711, -32'd5356, -32'd6902},
{-32'd8563, 32'd10975, 32'd2270, 32'd8537},
{-32'd3763, -32'd12700, -32'd6888, 32'd8194},
{32'd3558, -32'd73, 32'd843, -32'd1442},
{32'd5013, 32'd1088, -32'd8504, 32'd191},
{32'd8883, -32'd4168, -32'd8532, -32'd2101},
{-32'd1394, -32'd11181, 32'd2601, -32'd2496},
{-32'd2393, -32'd2058, 32'd3279, 32'd5857},
{32'd4019, 32'd13946, 32'd6607, 32'd5634},
{32'd2673, -32'd13891, -32'd15002, 32'd11237},
{32'd1115, 32'd2877, 32'd1962, -32'd7795},
{-32'd1715, -32'd1666, 32'd6248, -32'd4843},
{-32'd2647, -32'd6762, -32'd7959, 32'd658},
{-32'd5604, -32'd925, 32'd6961, 32'd14403},
{32'd9754, 32'd8450, -32'd863, -32'd2631},
{-32'd7703, -32'd2052, -32'd13444, 32'd81},
{32'd176, -32'd11219, 32'd1966, 32'd1559},
{-32'd5444, -32'd143, 32'd3641, -32'd2674},
{-32'd5336, 32'd4137, 32'd11241, -32'd9444},
{32'd10931, 32'd9404, 32'd24072, -32'd13958},
{-32'd256, -32'd6059, 32'd2447, -32'd3095},
{-32'd14303, -32'd2603, 32'd4517, -32'd7195},
{-32'd5732, -32'd4580, -32'd4954, 32'd9259},
{32'd1083, -32'd9205, 32'd12229, 32'd8959},
{-32'd2786, 32'd3067, 32'd2397, -32'd2073},
{32'd131, -32'd2509, -32'd1793, 32'd210},
{-32'd6242, -32'd3846, -32'd6783, -32'd3084},
{32'd7617, -32'd11432, -32'd3083, -32'd8668},
{-32'd3082, -32'd8518, -32'd5345, 32'd1664},
{32'd10590, 32'd5836, 32'd605, 32'd9085},
{-32'd1623, 32'd156, -32'd6322, -32'd6115},
{-32'd10641, -32'd9152, -32'd1790, -32'd10205},
{32'd1958, -32'd7536, -32'd1885, 32'd6305},
{32'd7579, -32'd328, -32'd1435, 32'd6066},
{32'd13700, -32'd3724, 32'd5837, 32'd11284},
{32'd6854, 32'd5003, 32'd6009, 32'd5049},
{32'd1852, -32'd1629, 32'd6187, 32'd637},
{32'd6092, -32'd2953, 32'd1555, 32'd622},
{32'd1143, 32'd5700, -32'd1424, -32'd1617},
{32'd10478, -32'd1235, 32'd1102, -32'd1646},
{-32'd5034, -32'd10379, -32'd1556, 32'd4074},
{32'd8411, 32'd9533, -32'd7954, 32'd5578},
{-32'd7659, 32'd1108, -32'd1182, -32'd5765},
{-32'd10745, 32'd4416, -32'd134, -32'd2794},
{32'd15012, 32'd3083, 32'd4979, -32'd4755},
{-32'd6650, 32'd4989, 32'd11722, -32'd6964},
{-32'd7010, -32'd726, 32'd2354, -32'd10293},
{-32'd13998, -32'd982, 32'd3263, 32'd4452},
{-32'd7335, -32'd3446, 32'd10944, -32'd3810},
{32'd630, -32'd3851, 32'd3038, 32'd3687},
{32'd16605, -32'd4266, -32'd5324, 32'd8280},
{32'd6513, -32'd1670, -32'd8337, 32'd12620},
{-32'd2180, -32'd1510, -32'd3020, -32'd2096}
},
{{32'd10208, 32'd5146, 32'd7575, -32'd2959},
{-32'd1042, -32'd3019, 32'd6807, -32'd2090},
{-32'd4263, 32'd3442, 32'd9893, 32'd7651},
{32'd2515, 32'd7400, 32'd4224, -32'd483},
{-32'd2671, 32'd1087, -32'd830, -32'd7473},
{-32'd4456, -32'd10238, 32'd5583, 32'd2137},
{32'd9984, -32'd3138, -32'd3443, -32'd1192},
{-32'd4153, 32'd195, 32'd8413, -32'd3131},
{32'd6409, -32'd440, 32'd6874, -32'd9106},
{32'd7886, 32'd8731, -32'd1069, 32'd1181},
{-32'd5865, 32'd3783, 32'd6168, -32'd3026},
{-32'd4212, 32'd4217, -32'd4061, 32'd3083},
{32'd349, -32'd7780, -32'd3190, -32'd71},
{32'd3797, 32'd4816, -32'd9209, 32'd219},
{-32'd7326, -32'd7610, 32'd267, -32'd2447},
{-32'd2658, -32'd13905, 32'd8551, 32'd7320},
{32'd6234, 32'd3296, 32'd3411, -32'd8367},
{-32'd403, 32'd603, -32'd342, 32'd8564},
{32'd2198, 32'd11355, -32'd9867, -32'd805},
{-32'd4789, 32'd5104, 32'd5027, -32'd3796},
{-32'd5047, 32'd6103, -32'd2702, -32'd1167},
{-32'd9650, 32'd1099, -32'd2587, 32'd3387},
{-32'd8827, 32'd5442, 32'd5682, -32'd36},
{32'd1512, 32'd6942, -32'd4741, -32'd8066},
{32'd1931, 32'd4100, 32'd1153, -32'd1576},
{32'd2033, 32'd7238, -32'd3237, 32'd3114},
{32'd3534, -32'd14163, 32'd9455, 32'd7827},
{-32'd4270, -32'd7326, -32'd4977, -32'd11530},
{32'd13651, 32'd11591, -32'd2056, -32'd247},
{-32'd5803, 32'd3559, -32'd15157, -32'd4380},
{32'd2179, -32'd8563, 32'd5263, -32'd6518},
{-32'd8018, 32'd3933, -32'd4280, 32'd3788},
{-32'd2065, 32'd2980, 32'd7380, 32'd6679},
{-32'd4522, -32'd8678, -32'd8099, -32'd3919},
{32'd4328, -32'd894, 32'd3745, -32'd3505},
{32'd6304, -32'd11647, 32'd2697, 32'd9294},
{-32'd6723, 32'd1403, -32'd949, -32'd1829},
{-32'd998, -32'd2000, -32'd8515, 32'd3700},
{32'd1440, -32'd1091, -32'd3354, -32'd11947},
{32'd4948, 32'd6286, 32'd4448, 32'd10560},
{32'd2624, 32'd11154, -32'd3848, -32'd547},
{32'd635, -32'd8702, 32'd980, 32'd3524},
{-32'd2756, -32'd1739, 32'd1088, 32'd432},
{-32'd3664, 32'd6460, 32'd333, 32'd689},
{32'd4506, 32'd4064, -32'd111, 32'd2479},
{-32'd4163, -32'd2238, -32'd3638, -32'd8506},
{-32'd8123, -32'd3150, -32'd10561, -32'd441},
{32'd375, -32'd7738, -32'd8116, 32'd1050},
{32'd16081, -32'd684, 32'd6940, -32'd10533},
{-32'd6966, -32'd12833, 32'd803, 32'd5574},
{32'd4407, -32'd1401, -32'd9808, -32'd9946},
{32'd9161, -32'd2457, -32'd8816, -32'd9040},
{-32'd2966, 32'd4253, -32'd9492, -32'd53},
{32'd9734, 32'd5073, 32'd3117, 32'd2787},
{32'd15148, -32'd531, 32'd5994, -32'd3143},
{-32'd5803, 32'd364, 32'd1294, -32'd6673},
{-32'd594, 32'd5650, 32'd1924, -32'd12145},
{-32'd6531, -32'd2357, -32'd8753, 32'd3221},
{32'd3951, -32'd181, 32'd6452, -32'd2845},
{-32'd2220, -32'd3365, 32'd2093, -32'd4021},
{32'd2378, -32'd5451, -32'd4070, -32'd4926},
{32'd6424, 32'd3082, 32'd5045, -32'd7473},
{-32'd1888, -32'd8494, -32'd4516, -32'd1673},
{-32'd5632, 32'd2629, 32'd759, 32'd6869},
{32'd1914, -32'd1691, -32'd2013, -32'd10016},
{32'd5160, -32'd5630, -32'd309, -32'd748},
{-32'd9611, -32'd6288, -32'd5301, 32'd3104},
{-32'd3657, -32'd1222, 32'd7052, -32'd4601},
{32'd5787, -32'd7750, -32'd9554, 32'd3597},
{32'd6369, -32'd6497, 32'd15789, 32'd1991},
{-32'd2523, 32'd12904, -32'd6244, -32'd9422},
{-32'd6858, -32'd6448, 32'd6115, 32'd4588},
{-32'd8628, -32'd477, -32'd3715, 32'd6992},
{32'd29, 32'd7597, 32'd5108, 32'd4554},
{32'd9800, 32'd8246, 32'd6107, 32'd2571},
{32'd12082, -32'd1214, 32'd1407, -32'd5143},
{-32'd1385, 32'd87, -32'd2174, 32'd1624},
{-32'd8383, -32'd9678, -32'd11069, -32'd10495},
{-32'd617, 32'd4017, -32'd9477, -32'd5688},
{32'd32, -32'd6584, 32'd9714, 32'd9524},
{32'd8516, -32'd8553, 32'd3811, 32'd1412},
{32'd3204, -32'd4369, -32'd13376, 32'd1716},
{-32'd13041, 32'd9331, 32'd3667, 32'd12212},
{-32'd2463, -32'd948, 32'd10250, 32'd6060},
{32'd9196, -32'd5379, 32'd2544, 32'd3656},
{32'd9758, 32'd402, 32'd5442, 32'd607},
{-32'd3109, 32'd2170, -32'd1871, -32'd5469},
{-32'd3581, -32'd8999, 32'd4348, -32'd1417},
{-32'd10153, 32'd240, -32'd4793, -32'd287},
{-32'd113, -32'd1138, -32'd11615, 32'd965},
{-32'd1981, 32'd301, -32'd4174, 32'd213},
{-32'd11178, -32'd7572, 32'd6209, 32'd7350},
{32'd2486, -32'd85, 32'd3047, -32'd1780},
{-32'd10227, 32'd6314, 32'd11279, -32'd581},
{-32'd5860, -32'd6509, 32'd4340, 32'd9246},
{32'd1784, 32'd6580, 32'd4619, -32'd4106},
{-32'd1104, -32'd783, -32'd1810, 32'd3231},
{32'd9763, 32'd10599, 32'd11157, 32'd4498},
{32'd5315, -32'd1451, 32'd1172, 32'd2040},
{32'd10050, -32'd3016, -32'd5246, -32'd3452},
{32'd2091, 32'd7425, -32'd997, -32'd624},
{32'd1323, -32'd16687, 32'd13869, 32'd957},
{32'd2619, 32'd13549, -32'd4133, -32'd2279},
{-32'd8683, 32'd4282, 32'd7102, -32'd4118},
{-32'd13092, -32'd2201, 32'd5055, -32'd4551},
{-32'd2073, -32'd8730, -32'd3817, -32'd1460},
{-32'd520, -32'd2689, 32'd3633, 32'd8989},
{32'd3812, -32'd2719, 32'd2179, -32'd1295},
{32'd671, 32'd8734, 32'd7301, -32'd288},
{32'd1815, -32'd3611, 32'd8940, -32'd589},
{32'd3328, 32'd8827, -32'd5824, -32'd3739},
{32'd5222, 32'd8893, 32'd2365, 32'd2063},
{32'd8578, 32'd6071, 32'd235, 32'd2428},
{-32'd1911, -32'd4363, -32'd2435, -32'd7748},
{-32'd11205, -32'd1426, 32'd12820, 32'd2564},
{32'd2770, -32'd5903, 32'd3749, 32'd1372},
{32'd3219, 32'd2939, 32'd6670, -32'd5413},
{-32'd2180, -32'd4318, -32'd2513, -32'd2275},
{-32'd2375, 32'd153, -32'd1016, -32'd8011},
{-32'd727, -32'd5625, 32'd5011, 32'd4644},
{32'd4917, 32'd3957, -32'd2770, -32'd3138},
{32'd7085, 32'd6054, 32'd3201, 32'd2175},
{32'd13779, -32'd2646, -32'd785, -32'd8893},
{-32'd5263, 32'd10134, -32'd875, 32'd4505},
{-32'd477, -32'd6750, -32'd1273, 32'd10024},
{32'd2124, 32'd3619, 32'd2618, -32'd1744},
{32'd10949, -32'd6612, 32'd8479, 32'd2808},
{32'd3244, 32'd4619, -32'd2737, -32'd6359},
{-32'd10066, -32'd334, 32'd7658, 32'd11525},
{32'd1639, -32'd5795, 32'd4483, -32'd8036},
{32'd5294, -32'd8093, 32'd1526, 32'd11546},
{32'd3585, -32'd158, -32'd468, -32'd1298},
{-32'd12958, -32'd6090, 32'd947, -32'd2046},
{32'd3038, 32'd14002, 32'd8283, -32'd937},
{-32'd1230, 32'd4073, -32'd4985, -32'd5491},
{-32'd10814, -32'd10197, -32'd5145, 32'd10483},
{32'd2854, -32'd14, -32'd6921, 32'd8380},
{32'd3380, -32'd5462, 32'd439, 32'd8294},
{32'd8442, -32'd12287, 32'd2519, -32'd16093},
{-32'd1882, -32'd2050, 32'd11405, -32'd5556},
{32'd10332, -32'd7342, -32'd1416, -32'd1689},
{32'd395, 32'd6621, -32'd10828, -32'd1228},
{-32'd6698, -32'd391, -32'd14263, -32'd1534},
{32'd5468, 32'd6923, 32'd8603, 32'd2491},
{32'd3743, -32'd421, -32'd560, 32'd1398},
{32'd1905, -32'd1418, -32'd1, -32'd7004},
{-32'd12291, -32'd2936, 32'd4157, 32'd1525},
{-32'd10021, 32'd5287, -32'd8914, -32'd3489},
{32'd12465, -32'd13813, 32'd5592, -32'd3499},
{32'd401, -32'd5381, 32'd2188, 32'd1182},
{-32'd5772, -32'd2622, 32'd622, -32'd1920},
{32'd12958, 32'd8417, 32'd5213, 32'd6600},
{-32'd9219, 32'd357, 32'd6198, 32'd931},
{32'd6015, -32'd9431, 32'd8053, 32'd11021},
{-32'd5408, -32'd817, 32'd1167, -32'd276},
{32'd2765, 32'd5516, 32'd4972, 32'd6423},
{-32'd1169, 32'd3637, 32'd4227, 32'd6555},
{-32'd7112, -32'd2199, 32'd9929, -32'd58},
{-32'd7543, -32'd2869, -32'd3337, -32'd2079},
{32'd9830, -32'd4525, -32'd3902, -32'd2387},
{-32'd8410, -32'd5888, 32'd12920, -32'd4493},
{32'd12553, 32'd9228, -32'd5547, 32'd1103},
{32'd2205, -32'd62, -32'd4498, -32'd1248},
{32'd5440, 32'd11786, -32'd2094, -32'd3816},
{32'd4171, -32'd4370, 32'd2971, -32'd2962},
{-32'd10261, 32'd6191, -32'd2958, -32'd2788},
{-32'd1360, -32'd4801, 32'd4989, 32'd6875},
{-32'd3334, -32'd3703, 32'd5923, -32'd2798},
{-32'd3309, -32'd13136, -32'd13400, -32'd1258},
{32'd1594, -32'd14246, -32'd2774, -32'd3036},
{-32'd4855, -32'd416, 32'd592, 32'd10988},
{-32'd3142, -32'd13868, -32'd5232, 32'd3488},
{32'd6859, -32'd1357, 32'd1447, 32'd1112},
{-32'd4002, -32'd6567, -32'd9337, -32'd8697},
{-32'd5489, 32'd2170, -32'd10867, 32'd5486},
{-32'd1086, 32'd180, -32'd1052, 32'd6088},
{32'd1716, 32'd7890, 32'd5648, -32'd7027},
{-32'd1025, 32'd10599, -32'd3904, 32'd1148},
{32'd12436, 32'd4628, -32'd638, 32'd1531},
{-32'd2403, 32'd7057, -32'd1138, -32'd1850},
{32'd782, 32'd3304, -32'd4999, -32'd6092},
{32'd1209, -32'd4771, -32'd133, -32'd1142},
{-32'd6822, 32'd2605, 32'd3040, 32'd5835},
{32'd577, -32'd7354, 32'd7923, 32'd3117},
{-32'd10759, 32'd1630, 32'd10723, 32'd8854},
{-32'd3623, 32'd4386, -32'd1429, -32'd3592},
{-32'd2438, -32'd5377, 32'd1446, 32'd1419},
{32'd8092, -32'd3060, 32'd1262, -32'd2821},
{-32'd2167, 32'd7129, -32'd2501, -32'd4575},
{32'd3042, 32'd6197, -32'd7436, -32'd621},
{32'd11657, -32'd3787, -32'd2660, -32'd830},
{-32'd2700, -32'd1921, -32'd10000, 32'd2065},
{-32'd6328, 32'd5062, 32'd7021, 32'd3872},
{32'd7331, 32'd2497, 32'd4092, 32'd5548},
{-32'd986, -32'd1500, 32'd2049, -32'd3323},
{32'd7927, -32'd4625, 32'd3293, 32'd8735},
{-32'd7919, -32'd7855, -32'd1072, -32'd6041},
{32'd7922, 32'd5282, 32'd4005, -32'd6563},
{-32'd1080, 32'd2774, 32'd2792, 32'd2507},
{32'd336, -32'd6571, 32'd12875, 32'd690},
{-32'd6005, 32'd5962, -32'd1270, 32'd1289},
{-32'd3681, -32'd2058, -32'd226, 32'd12168},
{32'd13849, -32'd594, -32'd233, 32'd5276},
{32'd565, 32'd3608, 32'd2439, 32'd1172},
{32'd5947, -32'd1753, -32'd18308, -32'd616},
{-32'd1907, 32'd9710, -32'd9149, -32'd2973},
{-32'd4099, 32'd1316, -32'd3670, -32'd1957},
{32'd973, -32'd2435, 32'd6183, -32'd9779},
{-32'd7987, 32'd915, -32'd10261, 32'd6798},
{32'd7588, -32'd1912, 32'd6899, -32'd5776},
{32'd1081, -32'd2819, -32'd1445, -32'd3955},
{-32'd286, -32'd8396, 32'd1102, -32'd6202},
{32'd9515, -32'd2308, 32'd6065, 32'd1213},
{32'd4510, 32'd11717, -32'd804, -32'd8822},
{-32'd8169, 32'd119, -32'd9707, -32'd3615},
{32'd2973, 32'd2542, -32'd350, -32'd2201},
{-32'd4056, 32'd6242, -32'd816, -32'd4487},
{-32'd6436, 32'd3304, 32'd2492, -32'd2388},
{-32'd5437, -32'd2064, 32'd2149, -32'd5127},
{32'd5289, -32'd1734, -32'd6376, -32'd623},
{32'd1807, -32'd8089, -32'd8177, -32'd3585},
{32'd10646, 32'd3144, 32'd4968, -32'd2326},
{32'd4467, 32'd7452, 32'd7496, -32'd3584},
{32'd5956, 32'd2268, -32'd2643, 32'd93},
{-32'd7823, -32'd5898, 32'd8749, 32'd5134},
{32'd1768, -32'd1174, 32'd3537, 32'd7980},
{-32'd1953, -32'd3397, -32'd12441, -32'd1986},
{32'd2900, -32'd5284, -32'd4506, -32'd5381},
{32'd5473, 32'd4191, -32'd963, 32'd8051},
{32'd964, 32'd968, -32'd1358, -32'd165},
{-32'd4414, -32'd9056, 32'd8831, 32'd1291},
{32'd6281, 32'd3284, 32'd3215, -32'd1166},
{32'd2840, -32'd8027, 32'd2244, -32'd525},
{-32'd8767, -32'd7400, -32'd1644, -32'd1974},
{32'd3170, -32'd5435, -32'd6104, -32'd2162},
{-32'd1088, 32'd6413, -32'd15316, -32'd1160},
{-32'd5328, -32'd5829, 32'd6299, 32'd5591},
{-32'd2349, -32'd2103, -32'd895, 32'd2806},
{32'd2941, -32'd9080, -32'd1568, 32'd1669},
{-32'd1649, -32'd5461, -32'd2815, -32'd502},
{32'd5495, -32'd2374, 32'd2281, 32'd8751},
{32'd6122, -32'd11014, -32'd4729, -32'd12395},
{-32'd9046, -32'd2244, 32'd4995, -32'd1309},
{-32'd6102, -32'd2964, -32'd2627, 32'd8855},
{32'd8076, 32'd1680, 32'd4375, 32'd1461},
{-32'd10050, 32'd5555, -32'd5925, -32'd2032},
{32'd1953, -32'd14606, 32'd3001, 32'd9160},
{-32'd9462, -32'd347, 32'd5182, 32'd3457},
{32'd2999, 32'd5868, -32'd4904, 32'd1412},
{-32'd7214, -32'd5868, -32'd2495, -32'd9170},
{-32'd590, -32'd6723, -32'd2118, 32'd6783},
{32'd189, 32'd2386, -32'd1780, 32'd6057},
{32'd1956, -32'd1701, -32'd5748, -32'd11463},
{-32'd10159, 32'd6038, 32'd1770, -32'd5457},
{-32'd6554, 32'd361, -32'd64, 32'd5490},
{32'd2733, 32'd1529, 32'd2808, 32'd2283},
{32'd1426, 32'd12338, 32'd13768, 32'd6432},
{32'd14453, 32'd585, -32'd3649, -32'd2758},
{-32'd3375, 32'd106, 32'd5184, 32'd9166},
{32'd3655, -32'd315, -32'd4899, 32'd10749},
{32'd3204, 32'd5544, 32'd4558, -32'd8119},
{32'd2949, 32'd458, 32'd3084, 32'd4574},
{32'd3995, -32'd7338, -32'd2287, -32'd1167},
{32'd6718, -32'd7640, -32'd6644, 32'd10524},
{32'd10495, 32'd2203, 32'd2448, -32'd6935},
{-32'd5728, -32'd4436, -32'd2994, 32'd2247},
{-32'd679, -32'd1465, -32'd2185, 32'd5095},
{32'd3606, -32'd3355, -32'd91, -32'd728},
{32'd6326, -32'd4211, -32'd1516, -32'd225},
{-32'd4876, -32'd2000, -32'd5957, -32'd1199},
{32'd3278, 32'd2344, -32'd5491, -32'd4823},
{32'd7876, -32'd2178, 32'd3285, -32'd11946},
{32'd3073, 32'd7765, -32'd5296, -32'd7051},
{-32'd3525, -32'd3700, 32'd4989, 32'd432},
{-32'd4785, -32'd6591, 32'd1591, -32'd7581},
{32'd10061, -32'd2402, -32'd1302, 32'd6863},
{32'd10858, 32'd4185, -32'd1182, 32'd1827},
{32'd2819, -32'd8298, 32'd633, -32'd1439},
{-32'd5648, -32'd5618, -32'd1677, -32'd524},
{-32'd4342, -32'd5869, 32'd4756, -32'd875},
{32'd287, 32'd14143, 32'd4856, 32'd5426},
{32'd2867, 32'd6549, -32'd10212, -32'd6339},
{-32'd1959, -32'd6769, 32'd4023, 32'd6294},
{-32'd14580, 32'd3835, -32'd1251, 32'd4926},
{32'd9867, -32'd6880, -32'd846, -32'd5403},
{-32'd6471, -32'd898, -32'd8728, 32'd2765},
{32'd2346, 32'd4006, -32'd16577, -32'd8162},
{32'd1693, 32'd3967, 32'd6415, 32'd2934},
{-32'd7936, -32'd4874, -32'd2121, -32'd6752},
{32'd8086, 32'd10083, 32'd4765, -32'd2851},
{32'd6895, 32'd9061, 32'd3358, -32'd5199},
{-32'd1229, 32'd3523, 32'd3566, -32'd3755},
{32'd8918, 32'd4439, 32'd1119, 32'd3890},
{32'd8078, -32'd6946, 32'd3456, 32'd7685},
{32'd1533, -32'd7843, -32'd7435, 32'd9242},
{-32'd2529, -32'd8260, 32'd5465, -32'd5044},
{32'd11148, 32'd4852, 32'd3967, 32'd5130},
{32'd3547, 32'd4902, 32'd1513, 32'd103},
{32'd3184, 32'd12500, -32'd6914, -32'd6561},
{32'd1939, -32'd7888, 32'd2249, 32'd1157}
},
{{32'd10202, -32'd746, 32'd1809, -32'd5638},
{-32'd5262, -32'd9542, -32'd2907, 32'd14771},
{-32'd1177, -32'd2458, -32'd3342, 32'd3521},
{32'd5467, -32'd13208, 32'd2198, 32'd5846},
{-32'd2904, 32'd13953, 32'd4191, -32'd14869},
{-32'd6179, -32'd11681, -32'd4450, 32'd5732},
{32'd2812, 32'd8478, 32'd2912, -32'd534},
{-32'd18516, 32'd3271, -32'd2982, -32'd4850},
{-32'd5372, -32'd861, -32'd3177, -32'd9222},
{32'd13631, 32'd4421, 32'd7916, 32'd6625},
{-32'd6355, -32'd7912, -32'd4666, -32'd2454},
{-32'd3037, 32'd5630, 32'd2746, 32'd8632},
{-32'd9030, 32'd957, -32'd6951, 32'd4603},
{32'd804, -32'd7872, 32'd2971, 32'd698},
{-32'd5642, -32'd3303, 32'd2230, 32'd7640},
{-32'd710, -32'd5051, 32'd10762, -32'd1802},
{32'd1426, 32'd5961, 32'd4558, -32'd15834},
{32'd15598, -32'd4988, -32'd1605, 32'd3285},
{-32'd2309, 32'd12581, 32'd6642, -32'd1619},
{32'd3981, 32'd6966, -32'd2130, -32'd11004},
{32'd567, 32'd2032, 32'd2655, 32'd7065},
{-32'd5921, -32'd11330, -32'd7961, 32'd10060},
{-32'd6299, -32'd1499, 32'd4276, -32'd4873},
{32'd460, -32'd2102, -32'd9299, -32'd2613},
{32'd4226, 32'd5112, 32'd15510, 32'd6946},
{-32'd9251, -32'd3957, -32'd684, 32'd258},
{32'd1201, -32'd4782, 32'd3909, -32'd3111},
{32'd1965, -32'd3793, -32'd6194, 32'd5595},
{32'd7214, -32'd1304, 32'd1064, 32'd9990},
{32'd4290, 32'd11893, -32'd4858, 32'd2165},
{-32'd8309, 32'd4510, -32'd338, 32'd4103},
{-32'd7953, -32'd5024, -32'd7068, -32'd14731},
{32'd8727, 32'd6371, 32'd10643, 32'd261},
{32'd592, -32'd1352, 32'd6776, -32'd713},
{32'd7907, 32'd4796, 32'd2013, -32'd4069},
{-32'd10012, 32'd1592, 32'd964, -32'd8200},
{32'd3342, -32'd11, -32'd3029, -32'd2287},
{-32'd852, -32'd4844, -32'd1064, -32'd235},
{32'd2890, 32'd3725, 32'd7785, 32'd4844},
{32'd3347, 32'd7096, 32'd13853, -32'd8534},
{32'd1804, 32'd2553, 32'd8215, 32'd2629},
{32'd38, 32'd15011, 32'd4207, -32'd10730},
{32'd10501, 32'd8096, 32'd9783, -32'd14482},
{-32'd7353, -32'd4040, 32'd8637, 32'd3782},
{-32'd12980, 32'd1340, -32'd7399, -32'd14933},
{-32'd4784, 32'd1260, 32'd4520, -32'd2749},
{-32'd3671, -32'd8823, -32'd7999, 32'd2713},
{32'd157, -32'd6305, -32'd13032, -32'd1244},
{-32'd1877, 32'd2560, 32'd3464, 32'd2908},
{-32'd9810, -32'd1245, 32'd3733, 32'd5167},
{-32'd1595, -32'd2215, -32'd11980, 32'd1212},
{-32'd5001, 32'd5799, 32'd666, -32'd1074},
{32'd2927, -32'd10218, -32'd1809, 32'd1258},
{32'd6443, 32'd423, -32'd4117, -32'd5824},
{-32'd293, -32'd3622, 32'd15662, 32'd1566},
{-32'd6731, -32'd308, 32'd1073, 32'd4546},
{32'd9516, 32'd1238, 32'd7825, 32'd5341},
{-32'd2487, -32'd1862, -32'd18396, -32'd10962},
{-32'd6354, -32'd9762, -32'd4103, -32'd9648},
{-32'd1568, 32'd11352, 32'd4147, -32'd1651},
{-32'd4149, 32'd292, -32'd2868, -32'd5568},
{-32'd12859, -32'd4708, 32'd2344, 32'd1699},
{-32'd6959, -32'd2038, -32'd12006, -32'd6565},
{-32'd609, -32'd9371, 32'd2137, -32'd4401},
{-32'd2969, 32'd13057, 32'd2944, 32'd2156},
{-32'd2882, 32'd9200, 32'd3581, -32'd375},
{-32'd7869, 32'd4166, 32'd655, 32'd8841},
{-32'd1459, 32'd344, -32'd379, 32'd7439},
{32'd1446, -32'd5804, 32'd1203, 32'd15743},
{-32'd5389, -32'd1055, -32'd4326, -32'd4530},
{-32'd6576, -32'd3660, 32'd1990, -32'd2986},
{32'd5700, -32'd9137, 32'd4486, 32'd3761},
{-32'd518, -32'd2199, -32'd8362, -32'd7479},
{32'd2771, 32'd874, -32'd4476, -32'd3116},
{32'd4332, 32'd5227, -32'd3442, -32'd2702},
{32'd2064, 32'd3391, 32'd4481, -32'd6011},
{-32'd2922, -32'd3776, -32'd6454, 32'd5405},
{-32'd9069, -32'd2366, -32'd9328, -32'd9520},
{32'd4374, -32'd2790, 32'd5702, 32'd605},
{32'd1226, -32'd6447, -32'd3325, 32'd8186},
{32'd4143, -32'd9285, 32'd3873, -32'd13417},
{32'd846, 32'd9540, 32'd6606, 32'd1645},
{-32'd795, -32'd7766, -32'd5817, 32'd1039},
{32'd2651, 32'd3196, -32'd3790, -32'd18039},
{-32'd6094, 32'd5558, 32'd8727, 32'd14900},
{-32'd839, 32'd10128, 32'd6553, 32'd685},
{-32'd257, 32'd10369, -32'd2706, 32'd266},
{-32'd12158, -32'd4469, -32'd5090, -32'd4013},
{32'd4232, 32'd2216, -32'd15167, -32'd4408},
{-32'd4828, 32'd2102, -32'd6513, -32'd11986},
{32'd6784, -32'd4554, 32'd4383, 32'd490},
{-32'd2695, 32'd5794, 32'd4523, -32'd4538},
{-32'd4350, -32'd2192, 32'd284, 32'd2457},
{32'd6220, 32'd6409, -32'd844, 32'd5201},
{32'd3524, -32'd1587, -32'd5074, 32'd7994},
{-32'd723, 32'd6509, 32'd429, 32'd456},
{32'd8903, 32'd908, 32'd5284, -32'd3250},
{-32'd7729, 32'd693, 32'd213, -32'd1167},
{-32'd5739, 32'd1402, -32'd9717, 32'd41},
{32'd5081, -32'd5772, 32'd6859, -32'd2618},
{-32'd7606, 32'd2066, -32'd3753, -32'd278},
{32'd2235, -32'd2551, 32'd3773, -32'd11852},
{32'd1271, 32'd3794, -32'd1127, -32'd1687},
{32'd1061, -32'd6811, -32'd2595, -32'd1230},
{32'd1089, 32'd4641, 32'd2555, -32'd4545},
{-32'd4809, -32'd259, 32'd7098, -32'd10929},
{-32'd3268, -32'd6142, -32'd9471, -32'd9186},
{-32'd11528, -32'd2975, 32'd3162, -32'd3869},
{32'd1082, -32'd4932, 32'd3196, -32'd4079},
{-32'd1595, 32'd1244, -32'd8628, -32'd5817},
{32'd8964, -32'd1673, -32'd9224, -32'd7697},
{32'd7047, 32'd3690, 32'd6703, -32'd3948},
{32'd7412, 32'd5805, 32'd10692, -32'd1453},
{-32'd387, 32'd6003, 32'd9343, -32'd11585},
{-32'd683, -32'd11552, -32'd3058, -32'd6909},
{-32'd3650, 32'd4667, 32'd4397, -32'd10194},
{32'd6175, -32'd4182, -32'd2762, -32'd1115},
{-32'd2895, -32'd1079, -32'd2712, 32'd2423},
{32'd12709, -32'd9715, -32'd525, -32'd2871},
{32'd14701, 32'd15490, 32'd309, -32'd369},
{32'd5682, -32'd5311, 32'd7489, -32'd6650},
{-32'd178, 32'd2585, 32'd1516, 32'd3907},
{32'd6826, -32'd799, 32'd9024, 32'd8927},
{32'd4272, 32'd4038, -32'd9825, 32'd5290},
{-32'd7610, 32'd3400, -32'd7327, 32'd7547},
{32'd1339, -32'd8070, 32'd1752, 32'd5521},
{-32'd3572, -32'd3891, 32'd1764, -32'd1784},
{-32'd8442, 32'd10534, 32'd446, -32'd1258},
{-32'd8480, 32'd1545, -32'd3511, -32'd477},
{-32'd6592, 32'd688, -32'd4013, -32'd8664},
{32'd5474, -32'd3469, -32'd7839, -32'd12329},
{-32'd4755, -32'd5492, 32'd3874, -32'd2891},
{-32'd6147, -32'd6277, -32'd6408, -32'd6524},
{32'd7376, 32'd2245, 32'd11036, 32'd12015},
{32'd5643, -32'd3340, 32'd5936, 32'd9308},
{32'd6018, 32'd1783, -32'd1697, 32'd6271},
{32'd9130, 32'd8782, 32'd3442, 32'd7552},
{32'd2864, -32'd4160, -32'd4480, -32'd2007},
{32'd7866, -32'd3700, 32'd216, -32'd2690},
{-32'd12409, -32'd6629, -32'd1241, -32'd4194},
{32'd3830, -32'd993, -32'd5455, -32'd1923},
{-32'd13002, 32'd9083, -32'd6756, -32'd2197},
{32'd14917, -32'd3886, 32'd4040, -32'd2972},
{-32'd13476, -32'd6777, -32'd8510, -32'd4829},
{32'd9899, 32'd7856, 32'd1586, 32'd126},
{32'd9297, -32'd2769, 32'd1577, -32'd3986},
{-32'd533, 32'd3047, 32'd1966, -32'd8261},
{32'd7540, -32'd12922, 32'd5297, 32'd2430},
{32'd141, 32'd4025, 32'd4705, 32'd2642},
{-32'd13028, -32'd12437, -32'd8701, -32'd849},
{-32'd4572, -32'd1451, -32'd6219, -32'd5173},
{32'd4109, -32'd2764, 32'd3973, -32'd7075},
{-32'd6550, -32'd4534, 32'd333, -32'd10329},
{-32'd263, -32'd7683, -32'd3168, -32'd6221},
{-32'd15041, -32'd7580, -32'd12039, -32'd7582},
{32'd1211, 32'd14794, 32'd4625, -32'd9839},
{-32'd8238, 32'd10549, 32'd4091, -32'd4284},
{-32'd5728, -32'd5011, -32'd4038, 32'd11027},
{32'd1407, -32'd4518, -32'd2894, -32'd6080},
{32'd3903, 32'd5287, -32'd2632, -32'd1027},
{-32'd1297, -32'd16591, -32'd5072, -32'd15328},
{32'd163, 32'd9712, 32'd1069, 32'd1538},
{32'd2771, -32'd6434, -32'd7629, -32'd9807},
{32'd3490, 32'd2546, -32'd2536, 32'd8070},
{32'd5918, 32'd5839, 32'd5628, -32'd1190},
{-32'd949, -32'd6152, 32'd282, 32'd6706},
{-32'd11507, -32'd15348, -32'd7849, -32'd2241},
{32'd1124, 32'd2579, 32'd186, 32'd2340},
{32'd3204, 32'd3754, 32'd1686, 32'd2841},
{32'd832, 32'd12789, -32'd3651, 32'd188},
{-32'd7095, 32'd619, -32'd8404, 32'd7887},
{32'd5541, 32'd15486, 32'd5369, 32'd2600},
{32'd10116, 32'd7238, 32'd7817, -32'd3794},
{-32'd8918, 32'd6317, -32'd7460, -32'd8230},
{-32'd506, 32'd1330, -32'd962, 32'd11135},
{-32'd2284, 32'd2895, 32'd7283, 32'd10156},
{-32'd9973, -32'd2833, 32'd12097, 32'd20722},
{-32'd289, 32'd5004, -32'd841, 32'd7430},
{32'd5883, 32'd3738, 32'd1346, 32'd3488},
{32'd389, -32'd7623, -32'd6514, 32'd7680},
{-32'd6961, -32'd6192, -32'd576, -32'd16143},
{-32'd7206, -32'd3291, 32'd3387, -32'd19649},
{-32'd14398, 32'd8578, 32'd1565, 32'd14720},
{32'd1542, 32'd4733, -32'd25, -32'd5984},
{32'd6418, -32'd13313, 32'd444, 32'd6926},
{-32'd4082, 32'd272, 32'd6151, 32'd8849},
{32'd172, -32'd5276, -32'd3039, -32'd345},
{32'd4600, 32'd168, 32'd9366, 32'd7382},
{32'd1076, 32'd6753, 32'd160, -32'd5767},
{32'd1863, 32'd824, 32'd1109, -32'd14965},
{32'd10232, 32'd5732, -32'd592, -32'd2799},
{-32'd11311, -32'd9427, -32'd3601, -32'd6573},
{32'd6391, -32'd1721, 32'd4358, 32'd1512},
{-32'd1870, 32'd4788, 32'd865, 32'd1880},
{-32'd2741, 32'd2916, 32'd3024, -32'd12061},
{32'd2257, -32'd3169, -32'd608, -32'd3409},
{-32'd4659, 32'd753, -32'd1766, -32'd4280},
{32'd5832, -32'd493, 32'd11794, 32'd14807},
{-32'd4506, 32'd3953, -32'd12453, 32'd2248},
{32'd1630, 32'd4276, 32'd2776, -32'd5325},
{-32'd8517, -32'd4681, -32'd6183, 32'd2185},
{32'd6896, -32'd7565, -32'd1407, -32'd17587},
{32'd1346, -32'd3243, 32'd67, -32'd1142},
{32'd8105, -32'd7730, -32'd2866, 32'd987},
{-32'd964, 32'd793, 32'd5153, -32'd2378},
{-32'd6862, 32'd8878, -32'd8499, -32'd3806},
{32'd6639, -32'd6092, 32'd444, 32'd6130},
{-32'd365, 32'd286, 32'd2776, 32'd8344},
{-32'd4355, -32'd6389, -32'd15171, -32'd11413},
{32'd2617, 32'd5254, -32'd3567, -32'd3730},
{32'd135, 32'd8456, 32'd4731, 32'd12834},
{32'd10280, 32'd8729, 32'd2939, -32'd3711},
{-32'd9726, 32'd3382, -32'd3360, 32'd1033},
{-32'd41, -32'd4496, -32'd152, 32'd4580},
{-32'd1364, -32'd13109, 32'd4044, -32'd1674},
{32'd10952, -32'd1884, -32'd4426, 32'd9220},
{32'd4756, -32'd284, 32'd8454, -32'd5680},
{-32'd1599, -32'd20639, -32'd6187, 32'd11281},
{32'd5026, 32'd2688, -32'd168, -32'd5288},
{-32'd25, -32'd4691, -32'd8506, -32'd831},
{32'd3504, 32'd2790, -32'd10331, -32'd6306},
{32'd102, -32'd3091, 32'd4259, 32'd3788},
{-32'd5389, -32'd72, 32'd3800, -32'd3433},
{-32'd5495, -32'd8988, 32'd1990, 32'd5834},
{-32'd1569, 32'd3038, 32'd4078, -32'd5774},
{-32'd5575, 32'd6282, 32'd4450, -32'd7394},
{-32'd4254, -32'd9487, -32'd886, -32'd4837},
{-32'd6737, 32'd5249, 32'd3554, -32'd2287},
{32'd4765, -32'd2940, -32'd4831, -32'd2449},
{32'd10149, 32'd857, 32'd8171, -32'd1455},
{-32'd4987, -32'd3565, -32'd1946, -32'd6595},
{32'd5434, 32'd3954, 32'd7900, 32'd5360},
{-32'd4650, -32'd6715, -32'd3185, 32'd204},
{-32'd2830, 32'd598, -32'd5529, -32'd15761},
{-32'd1404, 32'd10355, -32'd1512, 32'd8546},
{32'd5731, -32'd5025, 32'd7085, -32'd8913},
{32'd8514, 32'd2997, 32'd5508, 32'd8884},
{-32'd1909, 32'd21, -32'd5082, 32'd17615},
{32'd11500, 32'd1507, 32'd7631, -32'd3105},
{32'd2718, -32'd4405, -32'd1645, -32'd10712},
{32'd6425, 32'd2785, 32'd6418, -32'd2331},
{-32'd5725, 32'd2089, -32'd6625, -32'd10386},
{-32'd7340, -32'd16472, -32'd7181, -32'd2694},
{32'd1808, 32'd10273, 32'd2215, 32'd1632},
{32'd6020, 32'd3159, 32'd10497, -32'd630},
{32'd10953, 32'd390, -32'd3436, 32'd14690},
{-32'd862, 32'd4763, -32'd8513, -32'd1008},
{32'd7052, -32'd6984, -32'd3639, 32'd5234},
{-32'd4798, 32'd140, -32'd1566, 32'd9337},
{32'd2220, 32'd5884, 32'd1537, 32'd6951},
{-32'd2523, -32'd4712, -32'd2021, 32'd1760},
{32'd3337, -32'd2361, 32'd2730, 32'd11736},
{32'd2794, -32'd1686, 32'd6138, -32'd6440},
{-32'd2237, -32'd7393, 32'd999, 32'd6208},
{-32'd2181, -32'd8291, -32'd4001, -32'd17757},
{32'd8041, 32'd2471, -32'd3512, -32'd1682},
{-32'd695, 32'd2348, 32'd54, 32'd6744},
{32'd7675, -32'd2442, 32'd3076, 32'd60},
{-32'd8884, 32'd6414, -32'd4085, -32'd6418},
{32'd11695, 32'd10074, 32'd4475, 32'd2364},
{32'd4863, 32'd779, -32'd6976, 32'd4896},
{32'd7684, 32'd3527, 32'd2391, -32'd1786},
{-32'd8345, 32'd9734, -32'd5228, -32'd8176},
{-32'd4908, 32'd38, -32'd1918, -32'd959},
{-32'd7783, 32'd5671, 32'd6879, -32'd5892},
{-32'd13684, -32'd3990, -32'd6699, 32'd482},
{32'd22341, -32'd4439, -32'd4224, 32'd16099},
{-32'd6280, 32'd1390, -32'd2697, 32'd9607},
{-32'd3123, 32'd1137, -32'd3928, -32'd614},
{32'd71, 32'd12614, -32'd12196, -32'd9404},
{32'd5833, -32'd2194, 32'd1645, 32'd11779},
{32'd851, -32'd6776, 32'd2786, 32'd9089},
{-32'd9589, -32'd225, -32'd12488, -32'd6258},
{-32'd2350, -32'd700, 32'd873, -32'd17717},
{32'd10509, -32'd9164, 32'd1938, 32'd5481},
{-32'd5370, -32'd3345, -32'd2712, -32'd6757},
{32'd14587, 32'd8123, 32'd9263, 32'd2414},
{32'd2635, 32'd5633, -32'd3531, -32'd425},
{-32'd9959, -32'd4346, -32'd7030, -32'd2477},
{-32'd16444, 32'd10116, 32'd232, -32'd1399},
{-32'd451, 32'd1857, 32'd3164, -32'd4042},
{32'd8524, -32'd2191, 32'd4981, -32'd2646},
{-32'd4657, -32'd7100, 32'd5559, -32'd8710},
{32'd342, 32'd9486, -32'd3252, 32'd15327},
{32'd1318, 32'd8703, 32'd8121, -32'd2691},
{-32'd18797, 32'd4491, -32'd5927, 32'd251},
{32'd18304, 32'd2723, -32'd418, 32'd2055},
{-32'd17731, 32'd4761, -32'd1857, -32'd5294},
{32'd6192, 32'd13400, -32'd5812, -32'd5943},
{32'd1214, 32'd4929, 32'd3946, -32'd2894},
{-32'd3041, 32'd455, -32'd37, 32'd3715},
{32'd13988, -32'd1380, 32'd13439, 32'd16677},
{-32'd5523, -32'd6585, 32'd1649, -32'd3131},
{-32'd7574, -32'd4921, -32'd653, -32'd7304},
{-32'd10206, -32'd3109, -32'd4785, 32'd5344},
{-32'd187, 32'd97, -32'd4224, -32'd3410},
{-32'd723, -32'd8271, 32'd2682, -32'd9685},
{32'd7346, 32'd2117, 32'd5455, 32'd3052},
{-32'd309, 32'd1366, 32'd9074, 32'd4920},
{32'd7421, -32'd6347, 32'd1819, -32'd5736}
},
{{-32'd7008, 32'd7231, 32'd2282, 32'd4183},
{-32'd2312, -32'd12333, 32'd2502, 32'd3643},
{-32'd3616, 32'd4533, 32'd5426, -32'd814},
{32'd3288, 32'd2444, -32'd2353, 32'd4150},
{32'd5454, 32'd4546, -32'd4092, -32'd1102},
{-32'd4519, 32'd1831, -32'd3186, 32'd3648},
{32'd3332, 32'd1291, 32'd2071, -32'd3973},
{-32'd6540, -32'd6294, -32'd49, 32'd4293},
{-32'd12176, 32'd101, 32'd13543, -32'd1194},
{32'd13144, 32'd5662, 32'd1991, -32'd3578},
{32'd2694, 32'd176, 32'd519, 32'd5431},
{32'd10449, 32'd9590, -32'd2601, -32'd713},
{-32'd13848, -32'd3522, -32'd9325, 32'd211},
{-32'd10708, -32'd1264, 32'd3377, 32'd1553},
{-32'd15847, -32'd6818, -32'd2899, -32'd5874},
{32'd137, 32'd11040, -32'd5445, 32'd2422},
{-32'd4515, 32'd7936, 32'd2285, -32'd7743},
{32'd7792, -32'd1318, -32'd3790, 32'd930},
{32'd1563, 32'd4605, 32'd6264, 32'd7885},
{32'd12773, 32'd10271, 32'd4956, -32'd804},
{-32'd4756, -32'd8490, 32'd10144, -32'd1806},
{-32'd11441, -32'd14728, -32'd4644, 32'd9435},
{32'd4704, -32'd1389, -32'd5630, -32'd3785},
{32'd4283, -32'd7101, -32'd920, 32'd9111},
{32'd1677, 32'd10638, 32'd6627, -32'd4710},
{-32'd2224, -32'd7215, -32'd2679, -32'd7898},
{-32'd2457, 32'd1080, 32'd3382, -32'd4640},
{32'd10260, 32'd5961, -32'd1437, -32'd10806},
{-32'd7797, -32'd2189, 32'd9284, 32'd193},
{-32'd3001, 32'd5618, -32'd436, 32'd3933},
{-32'd1296, -32'd2121, 32'd194, 32'd13546},
{-32'd7198, -32'd7609, 32'd1164, -32'd708},
{-32'd2796, 32'd12964, -32'd8564, 32'd114},
{-32'd4100, -32'd1823, -32'd5981, -32'd1249},
{32'd9840, 32'd4231, 32'd376, -32'd6369},
{-32'd4264, 32'd4499, 32'd4021, 32'd2150},
{32'd9163, -32'd3287, -32'd3877, -32'd7338},
{32'd3954, -32'd4817, -32'd4798, 32'd3544},
{32'd1481, 32'd5825, -32'd1150, -32'd11359},
{-32'd2059, 32'd10624, 32'd3940, -32'd82},
{32'd4463, -32'd7543, -32'd3177, 32'd3827},
{-32'd1835, 32'd15153, -32'd5272, 32'd4306},
{32'd8251, -32'd836, -32'd1813, -32'd5764},
{-32'd1002, -32'd2102, -32'd4021, 32'd1443},
{32'd755, 32'd2477, -32'd15884, 32'd5830},
{-32'd155, -32'd11021, -32'd3061, 32'd3275},
{-32'd4930, -32'd10226, -32'd10986, 32'd11949},
{-32'd463, -32'd363, -32'd4183, 32'd9024},
{-32'd12846, 32'd3901, 32'd3429, -32'd2224},
{-32'd8657, 32'd5821, 32'd1357, 32'd1210},
{32'd37, -32'd6228, 32'd4635, -32'd708},
{32'd3207, 32'd6639, 32'd1583, -32'd13202},
{-32'd4882, -32'd15039, 32'd4148, -32'd573},
{-32'd15409, -32'd818, 32'd204, 32'd8351},
{32'd4508, 32'd3313, -32'd10707, -32'd6225},
{-32'd3144, 32'd3986, -32'd1858, 32'd9684},
{32'd3394, 32'd15303, 32'd3519, 32'd5764},
{-32'd5679, -32'd3855, -32'd6868, 32'd680},
{32'd348, -32'd5546, 32'd5920, 32'd13034},
{32'd9738, 32'd6567, 32'd2463, 32'd4517},
{32'd557, -32'd14226, -32'd1104, 32'd3206},
{32'd10729, -32'd5412, 32'd7769, -32'd2885},
{-32'd4796, -32'd6581, -32'd1156, -32'd407},
{-32'd1548, -32'd13204, 32'd9183, 32'd4031},
{32'd12180, 32'd1400, -32'd3273, -32'd3128},
{-32'd8315, 32'd8966, -32'd5378, 32'd1720},
{-32'd1531, -32'd5228, 32'd5142, 32'd6124},
{32'd5641, -32'd2904, -32'd8293, -32'd8283},
{-32'd2719, -32'd10625, 32'd3252, 32'd9932},
{32'd4165, -32'd5926, 32'd4729, 32'd8324},
{-32'd2685, -32'd1325, -32'd1743, -32'd7683},
{32'd442, -32'd6806, -32'd12601, 32'd3936},
{-32'd15300, -32'd7969, 32'd5607, 32'd676},
{32'd2818, 32'd5593, 32'd2955, 32'd5593},
{32'd6219, 32'd2871, 32'd888, -32'd1120},
{32'd6472, -32'd2324, 32'd9873, 32'd14668},
{-32'd3212, 32'd2337, 32'd12442, 32'd8074},
{32'd720, 32'd5413, 32'd7782, 32'd8686},
{-32'd15025, -32'd4631, 32'd11758, -32'd3214},
{-32'd977, 32'd6321, -32'd914, 32'd4028},
{-32'd5545, -32'd8461, -32'd3354, -32'd7911},
{32'd5060, 32'd3992, 32'd8124, 32'd7889},
{32'd1671, 32'd8389, 32'd1979, 32'd11610},
{-32'd7677, 32'd4978, -32'd10881, -32'd2982},
{-32'd3938, -32'd3343, -32'd2922, 32'd5337},
{32'd4293, -32'd1601, -32'd1087, -32'd12487},
{32'd7897, -32'd10217, -32'd1240, -32'd13775},
{-32'd8469, -32'd5956, -32'd1182, 32'd6907},
{32'd5563, -32'd1225, -32'd3960, -32'd655},
{-32'd4145, -32'd5675, -32'd117, 32'd9043},
{32'd14183, 32'd6407, -32'd11390, -32'd14015},
{32'd3407, -32'd9906, 32'd4812, -32'd8462},
{32'd10594, 32'd1113, -32'd2781, 32'd2534},
{32'd5927, 32'd9989, -32'd7298, -32'd4333},
{32'd15168, -32'd4177, -32'd9600, -32'd9475},
{32'd1859, -32'd13999, 32'd3753, 32'd3153},
{32'd15991, -32'd1240, -32'd4881, 32'd2945},
{32'd1520, 32'd3270, -32'd9148, -32'd1151},
{32'd7237, 32'd647, 32'd2075, -32'd7627},
{32'd1146, 32'd7980, -32'd3574, -32'd7303},
{32'd6906, -32'd17817, -32'd6131, -32'd14147},
{-32'd5684, -32'd2846, 32'd1761, -32'd120},
{32'd3269, 32'd7719, -32'd4166, -32'd935},
{-32'd4120, -32'd6094, 32'd19750, 32'd7227},
{32'd4885, 32'd1604, 32'd5331, -32'd1073},
{32'd15350, -32'd3207, -32'd12651, -32'd4196},
{-32'd697, 32'd2046, -32'd1290, 32'd646},
{-32'd21997, 32'd3264, 32'd2976, 32'd1198},
{32'd4808, 32'd1881, -32'd1958, 32'd2795},
{-32'd9717, -32'd5577, 32'd4131, -32'd4099},
{-32'd382, -32'd2912, -32'd5420, 32'd1658},
{32'd11245, -32'd4112, 32'd7767, 32'd9159},
{32'd4507, 32'd7949, 32'd11045, -32'd3465},
{32'd9842, 32'd1591, -32'd1029, 32'd919},
{-32'd2531, -32'd3713, 32'd6047, 32'd236},
{-32'd11638, 32'd354, 32'd4973, -32'd4503},
{32'd13814, -32'd7722, -32'd6198, -32'd9854},
{-32'd3399, 32'd970, -32'd4139, -32'd203},
{-32'd2535, 32'd5675, -32'd1252, -32'd938},
{32'd8238, 32'd11047, 32'd2087, -32'd1109},
{-32'd8690, -32'd2414, 32'd4101, -32'd6300},
{32'd2197, -32'd2461, 32'd4097, 32'd5709},
{-32'd14155, -32'd12909, -32'd1780, -32'd1467},
{32'd6540, -32'd6699, 32'd2171, 32'd763},
{32'd10243, -32'd5434, 32'd1061, -32'd7118},
{32'd2251, -32'd6170, 32'd2894, -32'd2620},
{32'd7191, 32'd860, 32'd8590, 32'd5646},
{-32'd9329, 32'd3219, 32'd1237, 32'd3354},
{32'd6417, -32'd6645, -32'd1902, -32'd5009},
{32'd599, 32'd5895, 32'd1095, -32'd715},
{-32'd15641, 32'd10808, -32'd72, 32'd7618},
{-32'd21, 32'd16420, -32'd5751, -32'd135},
{-32'd5725, -32'd3505, 32'd1841, 32'd846},
{-32'd15902, 32'd5491, 32'd5959, -32'd84},
{-32'd1562, 32'd4797, 32'd870, -32'd11906},
{-32'd11991, 32'd6020, -32'd6598, 32'd7481},
{32'd2810, 32'd722, -32'd4599, 32'd11945},
{32'd1585, 32'd2020, -32'd708, 32'd1277},
{32'd11523, 32'd7394, -32'd1984, 32'd4691},
{-32'd1203, 32'd920, -32'd812, 32'd11685},
{-32'd11262, -32'd2052, 32'd3248, 32'd7111},
{-32'd7255, -32'd9609, 32'd3978, 32'd16322},
{-32'd9975, -32'd92, -32'd3282, -32'd5599},
{32'd677, -32'd5074, -32'd12667, -32'd4502},
{32'd7208, -32'd2157, 32'd1814, -32'd8805},
{32'd2128, 32'd11523, -32'd11647, -32'd9656},
{-32'd4093, 32'd2649, -32'd8274, -32'd6992},
{-32'd6255, -32'd8669, -32'd3920, 32'd19749},
{-32'd4426, 32'd2484, 32'd12611, -32'd5017},
{-32'd12947, -32'd13807, 32'd4687, 32'd6292},
{-32'd717, 32'd11573, -32'd9545, -32'd2677},
{-32'd3730, 32'd9198, -32'd1524, 32'd5411},
{-32'd9678, 32'd10768, -32'd7189, -32'd5281},
{32'd2229, -32'd5324, -32'd6896, 32'd528},
{-32'd1999, -32'd5642, -32'd3913, 32'd1763},
{-32'd84, 32'd3471, -32'd8521, -32'd11817},
{-32'd201, 32'd9437, 32'd8400, -32'd3502},
{32'd10395, -32'd5613, -32'd1686, 32'd3083},
{32'd644, -32'd2034, -32'd12460, -32'd6877},
{-32'd6171, -32'd2914, -32'd3813, 32'd4134},
{-32'd4953, 32'd11819, 32'd3541, -32'd978},
{32'd4885, 32'd1244, -32'd5631, -32'd2824},
{32'd6683, -32'd3738, -32'd2391, -32'd214},
{32'd5747, 32'd7108, 32'd4815, -32'd3421},
{-32'd10818, 32'd340, 32'd3576, 32'd2234},
{32'd2059, -32'd7244, 32'd8753, -32'd333},
{-32'd7351, -32'd1760, -32'd7756, -32'd9867},
{-32'd3787, -32'd1344, 32'd3638, 32'd5168},
{-32'd5916, -32'd6334, -32'd5495, 32'd14347},
{-32'd1042, 32'd7231, 32'd2642, -32'd1662},
{-32'd5723, -32'd2739, 32'd9983, -32'd3318},
{-32'd2247, 32'd13267, 32'd6488, -32'd3014},
{32'd4613, 32'd5559, -32'd509, -32'd4833},
{-32'd6108, -32'd2685, 32'd9526, 32'd6179},
{-32'd2915, -32'd2745, -32'd442, 32'd4753},
{32'd12140, 32'd6994, -32'd5921, 32'd9966},
{-32'd1918, 32'd6380, 32'd5392, -32'd936},
{-32'd70, 32'd12542, -32'd151, 32'd732},
{-32'd4598, 32'd3348, 32'd470, 32'd4089},
{-32'd4129, -32'd1540, -32'd11334, 32'd3571},
{-32'd7258, -32'd1545, 32'd4182, 32'd10190},
{-32'd3533, 32'd5113, -32'd8276, -32'd317},
{-32'd4076, 32'd1572, 32'd8141, 32'd4226},
{-32'd2006, 32'd2759, -32'd3938, 32'd2014},
{-32'd4139, -32'd605, -32'd10044, 32'd4813},
{32'd7154, 32'd4501, -32'd10144, -32'd1865},
{-32'd3319, 32'd3781, 32'd1382, 32'd2548},
{32'd8248, 32'd11763, 32'd292, -32'd970},
{32'd7896, -32'd5922, 32'd7780, -32'd757},
{-32'd9446, -32'd264, -32'd5764, 32'd3229},
{-32'd13308, 32'd9741, -32'd3725, 32'd276},
{-32'd13496, -32'd3601, 32'd7979, 32'd4638},
{32'd3988, -32'd19661, 32'd4144, -32'd3738},
{-32'd4826, -32'd12396, 32'd1909, -32'd7935},
{32'd92, -32'd1117, -32'd6134, -32'd10944},
{-32'd42, 32'd4762, 32'd1136, -32'd4212},
{32'd3925, -32'd10835, 32'd1406, -32'd18244},
{32'd2836, 32'd5682, 32'd2489, -32'd3442},
{-32'd13169, 32'd9518, 32'd379, -32'd12149},
{32'd8409, 32'd8133, -32'd7651, 32'd1193},
{-32'd6388, -32'd8359, -32'd969, 32'd2995},
{-32'd4722, 32'd6645, 32'd2746, -32'd16366},
{32'd6811, 32'd4817, -32'd3581, 32'd7719},
{-32'd1935, 32'd2196, 32'd786, -32'd9094},
{-32'd5713, -32'd1966, 32'd7509, 32'd5755},
{32'd2317, 32'd5952, -32'd2379, -32'd9694},
{32'd6132, 32'd13034, 32'd1941, -32'd1482},
{-32'd3371, -32'd16052, 32'd1714, 32'd3658},
{32'd13823, -32'd6423, -32'd8737, 32'd2763},
{32'd2381, -32'd12199, -32'd10537, -32'd5112},
{32'd10881, 32'd19, -32'd8146, 32'd368},
{32'd17404, -32'd7896, -32'd3887, -32'd1518},
{-32'd5987, 32'd1442, 32'd2196, 32'd1842},
{-32'd3719, -32'd9577, 32'd10706, -32'd3759},
{32'd2265, 32'd10719, 32'd4487, 32'd2044},
{-32'd3992, -32'd12022, -32'd3373, -32'd7218},
{-32'd3703, 32'd8661, 32'd2985, -32'd6875},
{-32'd1164, -32'd1087, 32'd3286, 32'd6011},
{32'd8009, 32'd3602, 32'd2040, -32'd1269},
{-32'd3582, 32'd59, -32'd9584, 32'd4949},
{32'd1309, 32'd5159, -32'd13323, -32'd1492},
{32'd1949, 32'd2162, 32'd3732, 32'd3815},
{32'd3533, 32'd645, 32'd12474, -32'd5111},
{-32'd5937, -32'd2165, -32'd5720, 32'd3881},
{32'd1887, 32'd2776, 32'd1313, -32'd2373},
{32'd1293, 32'd4544, -32'd276, 32'd5107},
{-32'd4615, -32'd252, 32'd592, -32'd2443},
{-32'd654, -32'd9573, 32'd3572, -32'd2303},
{-32'd11579, -32'd1832, 32'd6505, 32'd6329},
{-32'd1694, 32'd2701, -32'd7438, 32'd1972},
{32'd944, 32'd3383, 32'd430, 32'd3111},
{32'd4922, 32'd2642, -32'd5018, -32'd2469},
{-32'd6411, 32'd257, 32'd2573, -32'd334},
{32'd5712, -32'd1061, -32'd16055, 32'd2490},
{-32'd2829, -32'd4208, -32'd9018, 32'd8432},
{-32'd4204, -32'd9925, -32'd5946, 32'd1765},
{32'd8187, 32'd2292, -32'd8714, -32'd2213},
{32'd609, -32'd2201, -32'd13884, -32'd12259},
{32'd1949, -32'd956, 32'd8075, 32'd7231},
{32'd2708, -32'd5500, 32'd1959, 32'd12518},
{-32'd4346, -32'd1593, -32'd199, 32'd804},
{32'd14268, -32'd5304, 32'd6342, 32'd11091},
{-32'd9459, -32'd16549, -32'd4047, -32'd527},
{-32'd3001, 32'd6481, 32'd4467, -32'd6767},
{32'd12454, 32'd6373, -32'd1602, 32'd1307},
{32'd205, 32'd2104, -32'd1936, 32'd1399},
{-32'd4181, 32'd12909, -32'd12978, 32'd3164},
{32'd5431, -32'd7811, 32'd1047, 32'd2345},
{32'd8194, -32'd1739, -32'd7512, 32'd6729},
{32'd7940, -32'd5180, -32'd6489, -32'd10643},
{32'd8101, 32'd4026, -32'd10577, -32'd3708},
{-32'd10320, -32'd10178, -32'd3324, -32'd9474},
{32'd11196, 32'd11872, -32'd10302, -32'd2083},
{-32'd13334, -32'd5308, -32'd4872, -32'd8072},
{-32'd8687, 32'd4272, -32'd6610, -32'd1826},
{-32'd2729, -32'd4181, 32'd3869, 32'd1258},
{32'd6415, -32'd897, 32'd1767, -32'd4304},
{32'd4549, 32'd2697, 32'd2662, 32'd3223},
{32'd2805, -32'd959, -32'd1972, 32'd11427},
{32'd6458, 32'd2011, -32'd3291, -32'd7174},
{-32'd7451, 32'd1953, -32'd1584, -32'd7887},
{32'd10583, -32'd5074, -32'd13610, -32'd4094},
{32'd3137, -32'd23491, 32'd6873, 32'd3091},
{32'd139, 32'd3422, 32'd28, 32'd8230},
{32'd9075, 32'd2049, -32'd4958, -32'd10114},
{32'd3206, 32'd11093, -32'd148, 32'd13955},
{32'd7765, 32'd6827, 32'd2901, 32'd4577},
{32'd5704, 32'd1197, 32'd1360, 32'd7724},
{-32'd12063, -32'd14079, -32'd4507, 32'd14362},
{32'd6300, 32'd6823, 32'd8441, 32'd6760},
{32'd9169, 32'd3230, 32'd10127, 32'd6740},
{32'd4642, 32'd6131, -32'd7874, -32'd333},
{-32'd2614, -32'd11695, -32'd7295, -32'd6005},
{-32'd8416, 32'd828, 32'd2509, -32'd2610},
{32'd6030, 32'd10399, 32'd3899, 32'd7558},
{32'd5980, 32'd1361, 32'd12433, 32'd6803},
{32'd8381, 32'd10096, 32'd1363, -32'd4300},
{-32'd5407, 32'd280, 32'd5911, -32'd4967},
{32'd867, -32'd12517, -32'd1589, 32'd9237},
{-32'd9778, -32'd7566, -32'd558, -32'd1352},
{32'd9121, -32'd4272, -32'd1497, -32'd3619},
{32'd1700, 32'd1445, 32'd12051, -32'd5670},
{32'd5306, 32'd5308, 32'd5575, 32'd220},
{-32'd11975, -32'd1982, 32'd11274, -32'd9946},
{32'd3400, 32'd18156, -32'd7368, -32'd6747},
{-32'd3827, -32'd6072, 32'd5906, 32'd5289},
{32'd3937, 32'd3182, 32'd7722, 32'd6438},
{-32'd1032, -32'd9335, -32'd12351, -32'd2944},
{32'd4161, -32'd4921, -32'd4240, -32'd9441},
{32'd1620, -32'd7210, -32'd1528, 32'd1969},
{32'd1572, 32'd40, 32'd515, 32'd6518},
{32'd11172, 32'd7458, 32'd9413, 32'd1313},
{-32'd15795, -32'd4656, 32'd7088, -32'd6596},
{32'd7412, -32'd13396, 32'd585, 32'd11126},
{-32'd10501, -32'd7296, -32'd4200, -32'd718},
{-32'd3972, 32'd6851, -32'd15105, -32'd9675},
{32'd8508, -32'd6128, -32'd3252, 32'd3472},
{-32'd1092, -32'd5719, 32'd8287, 32'd9971},
{-32'd3251, 32'd7041, 32'd11516, -32'd6565},
{-32'd262, 32'd3997, 32'd5862, 32'd11189}
},
{{32'd2063, 32'd2258, 32'd4771, 32'd1917},
{32'd7064, 32'd2035, -32'd5257, -32'd17467},
{32'd23219, -32'd1840, 32'd462, 32'd6487},
{32'd5754, 32'd8475, -32'd7902, 32'd2159},
{32'd9354, 32'd1755, -32'd4567, 32'd13192},
{32'd8582, -32'd5170, -32'd5017, -32'd11795},
{-32'd6338, 32'd2402, -32'd14028, 32'd9631},
{-32'd7889, -32'd8396, 32'd1001, -32'd4237},
{32'd2485, -32'd2691, -32'd2971, -32'd6051},
{32'd9331, 32'd4562, -32'd18, 32'd352},
{-32'd1738, -32'd5696, 32'd3908, -32'd1225},
{32'd5220, 32'd2382, -32'd14609, 32'd2232},
{32'd7011, -32'd15853, -32'd10971, -32'd564},
{-32'd6092, 32'd17077, -32'd9837, -32'd722},
{-32'd3275, -32'd4072, -32'd15211, -32'd2067},
{-32'd2205, 32'd5477, 32'd12771, -32'd15639},
{32'd11589, 32'd4035, 32'd5425, 32'd6837},
{-32'd13681, 32'd5756, 32'd11834, -32'd179},
{-32'd1897, 32'd12910, -32'd18066, -32'd684},
{-32'd7352, -32'd6078, 32'd12517, -32'd796},
{-32'd5376, -32'd2952, -32'd4007, 32'd1268},
{-32'd7790, -32'd6824, -32'd10427, -32'd2565},
{-32'd856, 32'd5628, 32'd328, 32'd1716},
{32'd593, -32'd840, 32'd9466, 32'd5990},
{32'd13486, -32'd945, 32'd3143, 32'd8116},
{32'd2714, 32'd3517, 32'd3880, 32'd6466},
{32'd793, -32'd130, 32'd3021, -32'd3074},
{32'd3911, -32'd6246, 32'd9302, -32'd1087},
{-32'd691, 32'd589, 32'd7603, -32'd12876},
{-32'd4888, 32'd2710, -32'd1114, -32'd1355},
{32'd9570, -32'd7359, -32'd14573, 32'd4415},
{-32'd3748, -32'd3883, 32'd1298, -32'd3187},
{32'd11728, -32'd3814, -32'd2110, 32'd3154},
{32'd2830, 32'd6525, 32'd2995, -32'd8312},
{32'd1093, 32'd3405, 32'd6896, 32'd7663},
{-32'd11934, -32'd8422, 32'd1469, -32'd2143},
{32'd6768, 32'd86, 32'd23128, -32'd10953},
{32'd6018, -32'd1815, -32'd6355, -32'd3875},
{32'd9759, 32'd7622, -32'd5295, 32'd2303},
{32'd7010, -32'd2904, -32'd2634, 32'd4676},
{-32'd5231, -32'd9050, 32'd6105, 32'd1073},
{32'd9899, 32'd11037, -32'd12585, 32'd949},
{32'd468, 32'd73, -32'd6639, 32'd6700},
{-32'd1949, 32'd11536, 32'd232, 32'd2487},
{-32'd3078, -32'd10658, 32'd15027, -32'd13006},
{-32'd1213, 32'd13808, -32'd10365, -32'd8245},
{-32'd17119, -32'd21178, -32'd4361, -32'd10281},
{32'd3220, 32'd6514, 32'd9060, 32'd1650},
{32'd5984, -32'd3072, 32'd2624, 32'd145},
{-32'd6224, 32'd3857, -32'd12803, -32'd3654},
{32'd8300, 32'd346, 32'd16, 32'd9741},
{32'd6318, 32'd2688, 32'd10099, -32'd547},
{32'd3902, 32'd1103, -32'd6724, 32'd10146},
{-32'd1024, -32'd7688, 32'd16011, 32'd8086},
{32'd3637, -32'd1507, 32'd911, 32'd107},
{32'd8964, 32'd3987, 32'd8896, -32'd8347},
{32'd1645, 32'd15983, -32'd10348, 32'd1904},
{32'd93, -32'd7649, 32'd6990, -32'd14096},
{-32'd2492, 32'd840, -32'd3300, -32'd14568},
{-32'd9480, 32'd20124, -32'd2044, -32'd1072},
{-32'd834, -32'd2431, -32'd13519, 32'd8291},
{-32'd2418, -32'd955, -32'd2209, 32'd5218},
{-32'd7675, -32'd2136, 32'd6761, -32'd7836},
{-32'd8527, -32'd4566, -32'd3685, -32'd10658},
{32'd19, -32'd3168, 32'd1948, -32'd5996},
{-32'd10792, 32'd2124, -32'd7184, 32'd9874},
{32'd9746, 32'd6489, 32'd2819, 32'd3723},
{32'd7536, -32'd11979, 32'd14110, -32'd125},
{-32'd7884, 32'd942, -32'd1879, -32'd9926},
{32'd745, -32'd135, 32'd17391, -32'd11613},
{-32'd8745, -32'd4493, 32'd10116, -32'd17553},
{-32'd1245, 32'd4469, -32'd911, -32'd2974},
{32'd4920, -32'd617, -32'd508, -32'd3320},
{-32'd6671, -32'd2534, -32'd16607, -32'd14018},
{-32'd4488, 32'd3997, -32'd3675, 32'd6237},
{-32'd1095, 32'd10945, 32'd15885, 32'd8021},
{32'd842, 32'd484, -32'd11187, -32'd17463},
{-32'd8511, 32'd15496, -32'd14034, -32'd5981},
{-32'd3721, 32'd271, -32'd6504, -32'd1166},
{32'd7432, 32'd14827, 32'd6822, 32'd15288},
{32'd7287, 32'd86, 32'd2281, -32'd2163},
{32'd3074, 32'd5964, -32'd9394, -32'd2877},
{32'd12150, -32'd1125, -32'd1466, -32'd1637},
{32'd6911, 32'd8936, 32'd14481, 32'd4475},
{32'd8960, 32'd3529, -32'd7395, 32'd11545},
{32'd9147, 32'd5247, -32'd4038, -32'd7580},
{32'd197, -32'd8189, 32'd9385, 32'd11344},
{-32'd8321, -32'd7894, 32'd8640, -32'd9079},
{-32'd784, -32'd2395, -32'd991, -32'd5152},
{32'd3416, 32'd9759, -32'd92, 32'd1704},
{32'd18816, -32'd139, 32'd4096, 32'd3381},
{-32'd15082, -32'd2858, -32'd16127, -32'd7942},
{-32'd1293, 32'd886, 32'd1817, 32'd6680},
{-32'd8901, 32'd2509, 32'd7309, 32'd14907},
{32'd1995, -32'd4148, 32'd17828, 32'd4443},
{-32'd5662, -32'd17119, 32'd582, -32'd1447},
{32'd5669, 32'd2389, -32'd16850, 32'd14748},
{32'd9522, -32'd13941, 32'd16493, 32'd9017},
{-32'd4412, -32'd9257, 32'd5023, -32'd7983},
{-32'd2337, 32'd6633, -32'd5697, 32'd9827},
{32'd1357, -32'd5614, -32'd7478, -32'd3889},
{32'd3408, -32'd1090, -32'd607, -32'd10554},
{32'd7847, 32'd3826, 32'd10287, -32'd1814},
{-32'd225, 32'd17727, -32'd5317, 32'd7581},
{-32'd11522, -32'd4400, -32'd10080, -32'd2662},
{-32'd18059, -32'd6247, -32'd10611, 32'd2327},
{-32'd2780, -32'd9060, 32'd6281, -32'd5970},
{-32'd7582, 32'd8257, 32'd3145, 32'd9058},
{32'd4435, 32'd13367, -32'd9626, -32'd1882},
{-32'd2351, -32'd7249, -32'd6420, -32'd3032},
{-32'd6310, 32'd8316, 32'd15659, 32'd1523},
{32'd1366, 32'd15980, 32'd11168, -32'd13677},
{32'd6058, 32'd9511, -32'd12128, 32'd13845},
{32'd1146, 32'd7664, -32'd8718, 32'd1689},
{32'd1314, -32'd5337, 32'd4545, 32'd3407},
{-32'd8929, -32'd1257, 32'd3814, -32'd5456},
{32'd6843, -32'd1095, 32'd4197, 32'd10639},
{32'd6617, 32'd1135, -32'd5876, -32'd2328},
{32'd2182, 32'd6546, 32'd9176, -32'd8078},
{-32'd8426, -32'd8398, -32'd6339, 32'd10279},
{-32'd1330, -32'd3869, -32'd6143, 32'd12731},
{32'd1903, 32'd7787, -32'd18217, 32'd13514},
{-32'd4386, 32'd3325, -32'd9167, 32'd3708},
{32'd2991, -32'd1448, 32'd14387, -32'd339},
{-32'd659, -32'd13652, -32'd17715, -32'd1840},
{32'd4645, -32'd8762, -32'd1812, 32'd521},
{32'd18939, -32'd744, 32'd2791, 32'd4107},
{-32'd11760, 32'd3676, -32'd1837, -32'd15030},
{-32'd416, 32'd4486, 32'd4153, -32'd4813},
{32'd11024, -32'd9793, 32'd3483, 32'd3060},
{-32'd11881, 32'd135, -32'd7538, 32'd16034},
{32'd7548, 32'd12360, 32'd11219, -32'd3128},
{-32'd11386, 32'd2627, 32'd6940, -32'd6985},
{32'd7710, -32'd1908, -32'd13222, -32'd853},
{32'd5466, -32'd13814, -32'd11648, -32'd8335},
{32'd9124, -32'd4100, 32'd2243, -32'd14886},
{-32'd1893, -32'd11132, -32'd2092, -32'd16384},
{32'd706, -32'd217, 32'd9618, 32'd4072},
{32'd10979, 32'd7815, -32'd6010, -32'd1653},
{-32'd7187, -32'd12840, 32'd16758, -32'd3510},
{-32'd16337, -32'd482, -32'd14885, -32'd7598},
{-32'd1253, -32'd6444, 32'd686, 32'd10798},
{-32'd2477, 32'd3163, -32'd2337, 32'd9600},
{-32'd10271, -32'd12295, 32'd7308, 32'd6028},
{32'd6599, 32'd4344, 32'd10043, 32'd6768},
{32'd6643, -32'd7958, 32'd10160, 32'd906},
{-32'd18329, -32'd3738, -32'd21472, 32'd9459},
{32'd239, 32'd1848, -32'd10810, 32'd1238},
{32'd5576, 32'd2424, 32'd7050, 32'd6770},
{32'd1925, -32'd3131, -32'd2376, 32'd3625},
{32'd1014, -32'd8292, 32'd13216, 32'd3691},
{-32'd5455, 32'd2576, -32'd10108, -32'd1420},
{-32'd3639, 32'd4000, -32'd12823, 32'd4489},
{32'd1724, 32'd4880, 32'd12956, 32'd4746},
{-32'd450, -32'd8378, 32'd3320, -32'd11978},
{32'd16111, 32'd5566, -32'd5257, -32'd7926},
{-32'd12399, -32'd3372, 32'd4388, -32'd3655},
{-32'd8497, 32'd6925, 32'd11801, 32'd3249},
{-32'd12123, -32'd3535, -32'd9589, -32'd1316},
{-32'd4188, -32'd2702, -32'd6272, -32'd13743},
{-32'd3299, 32'd2528, 32'd1583, -32'd1080},
{32'd7869, -32'd2703, 32'd13973, 32'd3088},
{-32'd2389, -32'd3454, 32'd8154, 32'd14172},
{32'd4517, -32'd3343, -32'd15288, -32'd58},
{-32'd10825, 32'd2935, -32'd3096, -32'd11148},
{-32'd9019, -32'd680, 32'd2439, -32'd1246},
{32'd7945, -32'd10767, 32'd10238, -32'd773},
{-32'd2561, -32'd2918, 32'd536, -32'd6917},
{32'd8975, -32'd3394, 32'd4898, -32'd1643},
{-32'd1243, -32'd2268, -32'd831, 32'd2309},
{-32'd535, -32'd8806, 32'd12910, 32'd975},
{32'd385, -32'd1755, 32'd17354, -32'd5118},
{32'd2919, 32'd7893, 32'd2648, -32'd3129},
{-32'd61, -32'd14306, -32'd12417, 32'd229},
{-32'd1843, -32'd6112, -32'd16629, 32'd7941},
{32'd938, 32'd2281, 32'd10401, -32'd5512},
{-32'd2669, 32'd8130, 32'd7555, -32'd2262},
{-32'd3851, 32'd2918, 32'd3368, 32'd6003},
{-32'd7570, 32'd8562, 32'd1844, -32'd811},
{32'd6813, -32'd9180, -32'd7804, 32'd5552},
{32'd2946, -32'd2327, 32'd12600, -32'd8184},
{-32'd3133, -32'd5588, -32'd2359, -32'd6503},
{32'd9967, -32'd12104, -32'd9773, -32'd21066},
{32'd4957, -32'd7215, -32'd4647, -32'd9361},
{32'd13730, -32'd15740, 32'd985, -32'd2682},
{-32'd5215, 32'd169, -32'd2234, 32'd2262},
{32'd1781, 32'd640, -32'd10396, -32'd4324},
{-32'd3175, 32'd7106, -32'd5043, 32'd1204},
{-32'd16791, -32'd2765, 32'd3219, -32'd7895},
{32'd11035, 32'd1446, 32'd3800, -32'd7344},
{-32'd1450, -32'd12486, 32'd7923, 32'd945},
{-32'd6491, 32'd1701, -32'd4001, -32'd7557},
{32'd2436, 32'd6264, 32'd4618, -32'd11347},
{32'd4495, 32'd1540, 32'd5842, -32'd1333},
{32'd4234, 32'd2079, 32'd8876, -32'd10567},
{32'd474, -32'd3774, 32'd2830, 32'd15425},
{-32'd572, 32'd1712, -32'd4523, 32'd923},
{-32'd1412, 32'd6745, -32'd11729, 32'd10180},
{32'd10129, -32'd22484, 32'd20249, 32'd6650},
{32'd3021, -32'd7555, 32'd13988, 32'd608},
{-32'd2270, -32'd4944, 32'd663, -32'd16679},
{32'd12016, -32'd13665, 32'd1282, -32'd750},
{-32'd11807, -32'd12015, 32'd6162, -32'd2221},
{32'd308, 32'd8003, -32'd10498, 32'd8741},
{-32'd17079, -32'd4867, -32'd1908, -32'd13099},
{32'd4672, 32'd9596, 32'd2895, -32'd2807},
{32'd1997, -32'd3472, -32'd12822, -32'd5997},
{32'd5123, -32'd7637, 32'd7875, -32'd6406},
{32'd2440, -32'd4606, 32'd6625, 32'd6970},
{-32'd930, -32'd3027, -32'd337, 32'd10432},
{-32'd1454, -32'd10737, 32'd6164, -32'd3133},
{-32'd1350, -32'd6568, 32'd16249, -32'd270},
{32'd1455, -32'd10098, 32'd2019, 32'd8194},
{-32'd11307, -32'd176, 32'd749, -32'd8961},
{32'd3199, -32'd2651, -32'd4696, 32'd920},
{32'd2746, -32'd9938, 32'd1242, -32'd2333},
{32'd3253, -32'd11316, 32'd15103, 32'd1020},
{-32'd3736, -32'd7209, -32'd7276, 32'd10416},
{-32'd3405, -32'd4256, -32'd8004, 32'd10656},
{-32'd14349, -32'd7545, 32'd6559, 32'd13259},
{-32'd5581, -32'd2453, -32'd1725, -32'd5317},
{-32'd4522, 32'd5590, 32'd485, 32'd8846},
{32'd7157, -32'd1668, -32'd1087, 32'd5908},
{32'd15231, 32'd5228, 32'd3449, 32'd8382},
{-32'd10640, -32'd5805, -32'd12371, 32'd401},
{-32'd7337, 32'd3242, 32'd952, 32'd9773},
{32'd14266, 32'd7754, 32'd4767, -32'd5630},
{32'd4476, 32'd1984, -32'd5837, 32'd2462},
{-32'd527, -32'd5109, 32'd9291, 32'd5146},
{32'd8906, -32'd6929, -32'd4045, 32'd5173},
{-32'd15152, -32'd9491, -32'd1132, -32'd17052},
{32'd13760, 32'd12133, -32'd10431, 32'd13927},
{-32'd6934, -32'd2695, -32'd2460, 32'd11379},
{32'd5597, -32'd9228, 32'd743, -32'd6550},
{32'd4997, 32'd1227, 32'd6737, -32'd10465},
{-32'd0, 32'd5351, -32'd6731, 32'd8233},
{-32'd7682, 32'd4558, -32'd961, -32'd5572},
{-32'd54, -32'd19760, -32'd8064, 32'd3323},
{32'd18712, 32'd17727, -32'd15631, 32'd3195},
{-32'd1751, 32'd1598, 32'd4577, -32'd1753},
{-32'd2913, -32'd3686, -32'd14627, -32'd7598},
{-32'd8493, -32'd6609, 32'd6803, 32'd130},
{32'd2933, -32'd1387, 32'd3595, 32'd721},
{-32'd1884, -32'd5557, 32'd4157, 32'd2790},
{32'd4180, 32'd7275, 32'd1171, -32'd7338},
{32'd7009, 32'd9700, -32'd18540, 32'd791},
{32'd11045, -32'd6026, 32'd14952, 32'd3643},
{-32'd9518, -32'd3796, 32'd8612, 32'd9173},
{-32'd3784, -32'd14147, 32'd9342, -32'd6071},
{-32'd15630, -32'd2805, -32'd6817, 32'd16250},
{32'd8244, -32'd3977, 32'd422, -32'd16628},
{32'd18143, 32'd3319, -32'd5880, -32'd7241},
{32'd7981, 32'd3534, 32'd18903, 32'd6147},
{-32'd11226, -32'd1484, -32'd8902, 32'd9862},
{-32'd15755, 32'd4357, 32'd3234, -32'd1106},
{32'd3825, 32'd8018, 32'd25184, -32'd12348},
{32'd2427, -32'd6233, 32'd7239, -32'd708},
{32'd8846, 32'd14534, -32'd1522, 32'd4776},
{-32'd8794, 32'd614, -32'd9338, -32'd12047},
{32'd2081, 32'd6151, 32'd5492, 32'd1125},
{32'd9731, -32'd3437, 32'd30830, 32'd9723},
{32'd7592, 32'd11108, 32'd16305, -32'd189},
{-32'd10145, -32'd1433, 32'd665, 32'd13570},
{32'd8736, -32'd2693, 32'd11577, -32'd14664},
{-32'd4787, -32'd4881, 32'd5697, -32'd5483},
{32'd7930, -32'd2688, 32'd6388, -32'd8238},
{32'd13276, 32'd8688, -32'd10189, -32'd3490},
{-32'd6201, -32'd611, -32'd6513, -32'd4346},
{-32'd14914, -32'd3073, 32'd8588, -32'd2480},
{-32'd5004, -32'd4765, 32'd11919, 32'd2441},
{32'd5261, 32'd2762, -32'd1884, -32'd3700},
{32'd2319, 32'd7627, -32'd2404, 32'd9304},
{-32'd6066, -32'd4318, 32'd7305, -32'd5266},
{-32'd3213, 32'd747, 32'd3495, 32'd20969},
{-32'd7269, 32'd4800, -32'd9962, 32'd2925},
{-32'd6395, -32'd8093, -32'd8081, -32'd2627},
{32'd9533, 32'd5936, 32'd195, 32'd5376},
{-32'd3435, -32'd2508, 32'd3622, -32'd780},
{-32'd1659, 32'd6034, 32'd4374, -32'd2139},
{-32'd8793, 32'd1487, 32'd367, -32'd568},
{-32'd1279, 32'd3695, 32'd11357, 32'd6808},
{-32'd4931, -32'd4591, -32'd5562, 32'd2149},
{-32'd5256, 32'd7933, 32'd4994, -32'd4764},
{-32'd13087, 32'd7377, -32'd8681, 32'd11150},
{-32'd1801, 32'd4455, 32'd14783, 32'd15016},
{32'd86, -32'd7355, 32'd6549, -32'd13322},
{32'd1085, 32'd13429, -32'd4745, -32'd7987},
{-32'd12257, -32'd12961, 32'd8275, -32'd3566},
{-32'd4588, -32'd1395, 32'd707, 32'd20495},
{-32'd7425, 32'd6857, -32'd2852, -32'd4706},
{-32'd2771, -32'd6377, -32'd16621, 32'd614},
{32'd1669, 32'd8259, -32'd4461, -32'd3482},
{32'd4174, 32'd7531, 32'd12621, 32'd5121},
{32'd5546, 32'd2052, -32'd3746, -32'd4726},
{32'd723, -32'd3210, 32'd12223, 32'd1420},
{32'd6850, -32'd3775, 32'd17865, 32'd7792},
{32'd4842, -32'd3383, 32'd11289, -32'd5884},
{32'd4918, -32'd3926, 32'd10079, -32'd759},
{32'd1162, 32'd8225, -32'd4851, -32'd5301},
{-32'd12974, 32'd2111, -32'd4433, -32'd6982}
},
{{32'd4705, 32'd4983, 32'd5130, 32'd867},
{-32'd5860, -32'd10239, 32'd3075, 32'd2644},
{-32'd8158, -32'd7588, -32'd7997, -32'd6675},
{-32'd130, 32'd8099, 32'd9221, 32'd2088},
{32'd10287, -32'd7692, 32'd799, 32'd4608},
{-32'd9720, 32'd2091, -32'd1454, 32'd10157},
{-32'd3505, 32'd5482, 32'd2152, 32'd5100},
{-32'd8173, 32'd3871, 32'd6277, 32'd2035},
{-32'd1155, -32'd6655, -32'd1948, 32'd5109},
{32'd11313, 32'd10452, 32'd1395, 32'd2907},
{-32'd13698, -32'd8004, -32'd7670, -32'd2225},
{32'd12406, 32'd2560, 32'd2674, -32'd3392},
{32'd7082, -32'd2227, -32'd611, 32'd10991},
{-32'd4886, -32'd4836, -32'd5741, -32'd4310},
{-32'd841, 32'd4073, -32'd3457, 32'd2216},
{-32'd21786, -32'd25905, -32'd2868, -32'd4418},
{32'd8545, 32'd4116, 32'd6989, 32'd1798},
{-32'd2103, 32'd10454, -32'd7506, -32'd6598},
{32'd632, -32'd1515, -32'd3006, -32'd741},
{-32'd13483, 32'd4039, 32'd7370, 32'd2714},
{32'd1790, 32'd4261, 32'd7638, -32'd4544},
{-32'd2679, -32'd1599, -32'd3115, 32'd6063},
{-32'd3035, -32'd5771, 32'd193, -32'd404},
{-32'd686, 32'd1696, -32'd9529, -32'd3039},
{32'd7992, 32'd7004, -32'd514, -32'd13},
{-32'd9375, 32'd9004, -32'd4178, 32'd4036},
{-32'd187, 32'd2724, -32'd3092, 32'd7674},
{32'd9645, 32'd3105, 32'd9303, 32'd1847},
{32'd7119, -32'd6894, -32'd1174, -32'd6947},
{-32'd11031, 32'd170, 32'd226, 32'd9653},
{32'd4765, -32'd5755, -32'd8445, 32'd8951},
{-32'd2589, -32'd1745, -32'd4558, 32'd7902},
{32'd14501, -32'd2714, 32'd1122, -32'd2045},
{-32'd1353, -32'd7486, 32'd559, 32'd3187},
{32'd8768, 32'd10577, 32'd7182, 32'd6909},
{-32'd4157, -32'd5339, -32'd3087, -32'd2345},
{-32'd5491, -32'd1028, 32'd79, -32'd1527},
{-32'd7378, -32'd7059, 32'd2010, -32'd2640},
{-32'd628, 32'd3252, 32'd11457, 32'd9570},
{32'd7734, 32'd13768, -32'd5659, 32'd4369},
{-32'd7879, 32'd4174, 32'd2170, 32'd225},
{-32'd2878, 32'd6002, -32'd5239, -32'd946},
{32'd3875, -32'd8273, 32'd3872, -32'd2121},
{-32'd6815, -32'd13080, -32'd765, 32'd6087},
{-32'd5976, 32'd6992, -32'd4764, 32'd4892},
{32'd1949, -32'd534, 32'd2807, 32'd5893},
{32'd703, 32'd4238, -32'd6150, -32'd5179},
{32'd1465, 32'd3165, -32'd6891, -32'd6769},
{32'd3646, 32'd4058, -32'd10707, -32'd1277},
{-32'd12565, -32'd6062, 32'd8106, -32'd1753},
{32'd7177, -32'd8778, -32'd10886, 32'd9054},
{32'd5531, 32'd9516, 32'd2247, -32'd373},
{32'd3154, -32'd13158, -32'd16547, -32'd17727},
{32'd3027, -32'd1593, -32'd5021, -32'd10099},
{-32'd244, -32'd2807, -32'd4892, -32'd431},
{-32'd3488, -32'd8154, 32'd5815, 32'd6780},
{32'd10512, 32'd703, 32'd2589, -32'd297},
{-32'd7215, -32'd11054, -32'd7508, 32'd3944},
{-32'd9270, 32'd1983, -32'd7701, -32'd5376},
{-32'd4147, 32'd8047, -32'd3353, 32'd10792},
{32'd1756, 32'd12427, -32'd453, -32'd819},
{-32'd4567, 32'd2405, 32'd2248, -32'd3210},
{-32'd11721, -32'd9489, -32'd4790, 32'd7419},
{-32'd4544, -32'd4201, -32'd375, 32'd8646},
{32'd4563, 32'd2808, -32'd7576, -32'd10186},
{32'd15081, 32'd11390, 32'd10296, 32'd211},
{32'd3622, 32'd10615, 32'd5594, 32'd12143},
{32'd1336, 32'd10845, 32'd418, 32'd2615},
{-32'd5644, -32'd2985, 32'd5869, -32'd4360},
{32'd1878, 32'd13018, -32'd4007, 32'd14153},
{32'd555, 32'd3345, 32'd2706, 32'd10494},
{-32'd11076, -32'd11278, 32'd7072, 32'd4695},
{-32'd18442, -32'd4502, -32'd9579, 32'd9157},
{-32'd5695, -32'd1669, 32'd9566, -32'd6003},
{32'd12186, 32'd10349, 32'd7516, 32'd1549},
{-32'd5223, -32'd3647, 32'd4460, 32'd5831},
{-32'd14234, -32'd3370, -32'd1347, -32'd5479},
{32'd10259, -32'd8764, -32'd7706, -32'd10052},
{32'd5110, 32'd6266, -32'd789, 32'd2456},
{32'd2321, -32'd559, -32'd1860, 32'd284},
{32'd268, 32'd139, 32'd5383, -32'd1553},
{-32'd3128, -32'd3468, -32'd5085, -32'd7493},
{32'd1782, -32'd8944, 32'd234, 32'd2338},
{-32'd11555, -32'd13963, 32'd9629, -32'd3088},
{32'd393, -32'd7217, 32'd5538, -32'd3196},
{32'd1664, -32'd1811, -32'd4986, 32'd21159},
{32'd10758, 32'd2163, -32'd6301, -32'd7603},
{-32'd13634, -32'd6838, -32'd1424, -32'd309},
{-32'd5126, -32'd8134, -32'd15077, -32'd1563},
{-32'd549, 32'd7942, -32'd4997, 32'd4850},
{-32'd13, 32'd8296, -32'd3629, -32'd7684},
{-32'd370, -32'd1684, -32'd4216, 32'd4149},
{32'd2768, 32'd12235, -32'd6654, -32'd22},
{32'd4439, -32'd240, 32'd4399, -32'd937},
{-32'd2317, -32'd2997, -32'd4520, -32'd3333},
{-32'd5232, -32'd1479, -32'd66, 32'd10161},
{32'd7596, 32'd6509, 32'd732, -32'd1819},
{-32'd8976, 32'd5362, -32'd12426, 32'd3869},
{32'd7880, 32'd7300, 32'd6735, -32'd1799},
{-32'd2875, 32'd2656, 32'd2265, 32'd4296},
{-32'd4930, -32'd6008, -32'd6489, -32'd5363},
{-32'd5829, -32'd9827, 32'd785, -32'd1939},
{32'd5324, 32'd7056, -32'd7684, -32'd3489},
{32'd8654, 32'd4363, 32'd12526, -32'd2834},
{32'd10520, 32'd958, 32'd9247, 32'd99},
{32'd10578, 32'd40, -32'd6154, -32'd904},
{-32'd5248, -32'd3287, -32'd7504, 32'd556},
{-32'd3454, -32'd7475, 32'd7607, -32'd1224},
{32'd2059, 32'd14658, -32'd732, 32'd4364},
{-32'd10189, -32'd14280, 32'd2175, 32'd5366},
{-32'd6289, 32'd571, 32'd8424, -32'd5317},
{-32'd3103, 32'd2994, 32'd6265, -32'd1421},
{32'd3066, 32'd5152, 32'd2407, 32'd2223},
{-32'd3643, 32'd7092, 32'd3058, 32'd5421},
{32'd3157, -32'd10569, -32'd3147, -32'd1344},
{-32'd5140, -32'd5840, 32'd9951, -32'd930},
{32'd1274, -32'd7935, 32'd7546, 32'd47},
{-32'd3658, 32'd4774, -32'd48, 32'd4667},
{32'd1397, -32'd7964, 32'd10546, 32'd1886},
{32'd11746, 32'd8607, 32'd1330, 32'd5060},
{32'd15608, 32'd1392, 32'd2831, -32'd3372},
{32'd5551, -32'd1491, -32'd1223, -32'd2607},
{32'd4372, 32'd539, 32'd16400, 32'd4363},
{32'd9288, -32'd1051, -32'd1957, 32'd4878},
{32'd3063, -32'd473, -32'd4130, -32'd13588},
{-32'd1435, 32'd1901, 32'd2596, 32'd6411},
{-32'd12149, -32'd2027, -32'd3151, 32'd4017},
{32'd4177, -32'd3001, 32'd13191, 32'd1758},
{-32'd2131, -32'd9897, -32'd1183, -32'd7735},
{32'd10041, 32'd6540, 32'd6072, -32'd4759},
{32'd3046, 32'd1555, 32'd8918, 32'd7659},
{-32'd6400, 32'd473, 32'd489, 32'd2606},
{-32'd7164, -32'd6523, -32'd98, 32'd2878},
{32'd2136, -32'd1882, -32'd2628, 32'd3796},
{32'd10538, -32'd725, -32'd172, 32'd9199},
{-32'd416, -32'd8428, -32'd4150, 32'd4330},
{32'd7116, 32'd4210, 32'd1834, 32'd16629},
{32'd9060, 32'd2100, 32'd5047, -32'd2116},
{32'd300, -32'd1597, -32'd1992, -32'd7903},
{-32'd3775, -32'd2025, 32'd408, 32'd1345},
{32'd1242, -32'd2777, 32'd4572, 32'd1903},
{-32'd1885, 32'd1622, -32'd5810, -32'd1741},
{32'd4255, -32'd6533, 32'd5771, -32'd4873},
{-32'd13289, -32'd2065, -32'd1793, -32'd7819},
{32'd8112, 32'd15643, -32'd2768, 32'd5969},
{32'd9985, 32'd5768, 32'd188, -32'd2833},
{32'd835, -32'd17724, -32'd7932, 32'd771},
{32'd6376, 32'd2244, 32'd2193, 32'd12517},
{-32'd1801, 32'd7559, 32'd767, 32'd2298},
{-32'd2892, -32'd3915, 32'd1617, 32'd3500},
{-32'd6959, -32'd1003, -32'd5106, -32'd6632},
{32'd5670, 32'd686, 32'd4714, -32'd6850},
{-32'd6634, -32'd13626, 32'd15581, -32'd4091},
{-32'd5998, -32'd8947, -32'd7236, -32'd10944},
{-32'd12798, 32'd3014, -32'd6951, -32'd1522},
{32'd9825, 32'd5994, 32'd2996, -32'd8393},
{32'd8772, 32'd1271, 32'd6207, -32'd4228},
{32'd1789, 32'd19793, 32'd4177, -32'd307},
{32'd4600, -32'd312, 32'd4857, -32'd7424},
{32'd27, 32'd3838, -32'd510, 32'd3060},
{32'd3776, -32'd9837, 32'd2235, -32'd3053},
{32'd12511, 32'd2451, -32'd10908, 32'd746},
{-32'd2057, -32'd8478, 32'd4968, 32'd314},
{32'd8757, 32'd7971, 32'd4004, -32'd4741},
{32'd7356, 32'd3602, -32'd1596, 32'd6497},
{-32'd7365, 32'd9598, 32'd2092, 32'd6314},
{32'd1549, 32'd6926, -32'd10325, -32'd2657},
{-32'd5433, -32'd3780, -32'd537, -32'd2972},
{-32'd5476, -32'd226, 32'd4524, -32'd7045},
{-32'd1084, -32'd7020, -32'd790, 32'd5665},
{-32'd7821, 32'd7813, -32'd6212, -32'd11222},
{32'd4793, 32'd12658, -32'd784, -32'd887},
{32'd6064, 32'd10272, 32'd8753, 32'd5601},
{32'd1915, 32'd2283, -32'd12834, -32'd980},
{32'd6844, 32'd5315, 32'd289, -32'd1964},
{-32'd5869, -32'd4571, -32'd5129, -32'd2256},
{32'd3826, 32'd11741, 32'd7209, 32'd859},
{32'd7778, 32'd1952, 32'd6129, 32'd8234},
{32'd985, -32'd604, 32'd5565, -32'd2379},
{-32'd5965, -32'd9694, -32'd8309, -32'd11471},
{-32'd4316, -32'd3391, 32'd1496, -32'd4862},
{-32'd4169, -32'd15859, -32'd3186, -32'd4480},
{32'd1395, -32'd5487, -32'd7445, -32'd1841},
{32'd7988, 32'd2911, 32'd5135, 32'd9711},
{-32'd6984, -32'd2682, -32'd6445, -32'd14619},
{32'd538, 32'd1424, 32'd11723, -32'd2942},
{32'd6560, 32'd13056, 32'd9475, 32'd9764},
{32'd11264, -32'd13803, 32'd4829, -32'd2318},
{-32'd3733, -32'd7729, -32'd1813, 32'd3754},
{32'd1768, -32'd46, 32'd415, 32'd1425},
{32'd10404, 32'd8740, -32'd7229, -32'd5470},
{32'd2264, -32'd6063, -32'd5018, 32'd4019},
{-32'd4449, -32'd3201, -32'd7913, 32'd324},
{32'd15588, 32'd1049, -32'd1251, 32'd2724},
{-32'd13112, -32'd5456, 32'd9991, 32'd10562},
{-32'd5116, 32'd9043, 32'd3494, -32'd4622},
{-32'd10122, 32'd1519, 32'd6408, -32'd5015},
{32'd15906, -32'd7114, 32'd10274, -32'd3430},
{32'd2152, 32'd5981, -32'd4556, -32'd7446},
{32'd428, 32'd7669, 32'd9223, -32'd1092},
{-32'd7860, -32'd10272, -32'd3276, -32'd5104},
{-32'd6557, 32'd10103, -32'd8099, 32'd17666},
{32'd805, -32'd4995, 32'd1825, 32'd389},
{32'd12756, 32'd4251, 32'd7274, 32'd3792},
{-32'd4824, -32'd4069, -32'd1106, 32'd365},
{32'd3900, 32'd4981, 32'd3507, 32'd4810},
{32'd657, -32'd1462, 32'd8462, -32'd7652},
{-32'd1604, -32'd6297, 32'd4325, -32'd6848},
{-32'd5958, 32'd1585, -32'd11262, -32'd1855},
{32'd4667, 32'd6283, 32'd1299, 32'd3004},
{-32'd7240, 32'd5569, 32'd2295, -32'd4553},
{-32'd4398, -32'd2475, 32'd1078, 32'd9750},
{-32'd1813, -32'd2481, 32'd3003, 32'd5638},
{-32'd3081, 32'd19331, 32'd2712, -32'd5788},
{-32'd3039, -32'd2895, -32'd8306, -32'd7758},
{32'd3273, -32'd1098, -32'd10010, -32'd1392},
{-32'd7333, 32'd13374, 32'd5415, 32'd8783},
{32'd1967, -32'd9072, 32'd613, -32'd3457},
{-32'd5272, 32'd9770, 32'd8593, 32'd13730},
{32'd4391, 32'd1078, 32'd9348, 32'd3413},
{32'd654, -32'd8232, 32'd2714, -32'd233},
{32'd13051, -32'd9359, -32'd556, -32'd7325},
{32'd10088, 32'd6818, 32'd3766, -32'd1163},
{32'd1639, -32'd4066, -32'd5900, -32'd8212},
{-32'd4649, -32'd12051, -32'd7723, -32'd909},
{-32'd11073, 32'd2052, -32'd4205, 32'd1456},
{32'd6497, -32'd8046, -32'd2254, -32'd7501},
{-32'd9381, -32'd6422, -32'd9508, 32'd2523},
{32'd6300, 32'd2051, 32'd9090, 32'd4664},
{32'd4420, -32'd2252, 32'd9978, 32'd6542},
{-32'd5204, 32'd3326, 32'd2343, 32'd10497},
{-32'd2581, -32'd1023, -32'd8652, -32'd4900},
{-32'd1013, -32'd4446, -32'd1174, -32'd1702},
{-32'd13376, -32'd5224, -32'd2910, -32'd7475},
{32'd3197, 32'd2296, -32'd3284, -32'd4551},
{-32'd8636, -32'd12399, -32'd7443, -32'd2280},
{32'd4519, -32'd9296, 32'd8744, -32'd13006},
{32'd8232, -32'd5369, -32'd9601, 32'd631},
{32'd3128, -32'd1385, 32'd9281, 32'd6520},
{-32'd16556, -32'd5358, -32'd7785, -32'd4603},
{32'd9392, -32'd3475, 32'd5077, 32'd740},
{-32'd12423, 32'd4921, -32'd2566, -32'd204},
{-32'd11823, -32'd13547, -32'd5117, 32'd2174},
{-32'd6347, -32'd6640, -32'd3110, -32'd5584},
{32'd8259, 32'd9258, 32'd11271, 32'd6335},
{32'd9236, 32'd10788, -32'd2802, -32'd4719},
{-32'd4653, -32'd5258, -32'd6622, -32'd9545},
{-32'd420, 32'd1299, -32'd5949, 32'd1453},
{-32'd7282, 32'd4444, -32'd9346, -32'd16494},
{-32'd8754, 32'd227, 32'd11403, 32'd5336},
{-32'd7712, -32'd11713, -32'd7759, -32'd8366},
{32'd18169, 32'd5883, -32'd5097, -32'd2172},
{32'd11458, 32'd2391, -32'd1231, 32'd5508},
{32'd5558, -32'd8593, -32'd1756, 32'd3478},
{-32'd10585, -32'd11112, 32'd5782, -32'd1645},
{32'd8780, 32'd14300, 32'd4911, 32'd11930},
{-32'd4941, 32'd10153, 32'd4112, 32'd313},
{32'd4336, 32'd358, 32'd3892, 32'd5825},
{-32'd4730, -32'd6303, -32'd5135, -32'd6325},
{-32'd940, 32'd1939, 32'd5888, 32'd7040},
{-32'd8371, 32'd4733, -32'd3770, -32'd3296},
{32'd8996, -32'd12807, 32'd1052, 32'd884},
{-32'd4461, -32'd4362, -32'd4692, -32'd10160},
{-32'd2702, 32'd5467, -32'd2694, -32'd6329},
{-32'd51, 32'd9337, 32'd3198, -32'd1855},
{-32'd5308, -32'd7822, -32'd4812, -32'd868},
{32'd3176, 32'd1301, 32'd2275, 32'd193},
{-32'd6000, 32'd4308, 32'd5460, -32'd886},
{-32'd14316, -32'd8687, -32'd4415, 32'd1045},
{-32'd963, -32'd3266, -32'd9710, -32'd892},
{32'd2978, 32'd11807, 32'd4516, -32'd3006},
{32'd8918, 32'd3794, 32'd6307, 32'd2918},
{-32'd4104, -32'd805, 32'd3419, 32'd1817},
{-32'd6417, -32'd10366, 32'd253, 32'd6431},
{-32'd2530, -32'd10660, 32'd8640, -32'd983},
{-32'd11241, -32'd3202, -32'd1128, 32'd228},
{32'd9932, 32'd11740, 32'd6270, 32'd4886},
{-32'd2076, -32'd2439, 32'd14296, -32'd4314},
{-32'd5958, -32'd9822, -32'd7436, -32'd5260},
{-32'd3583, -32'd6171, -32'd1802, 32'd7785},
{32'd16661, 32'd7755, -32'd6173, -32'd1568},
{-32'd4834, -32'd4602, -32'd30, 32'd6908},
{-32'd3229, -32'd7398, 32'd10707, -32'd6014},
{32'd6828, 32'd3590, -32'd1484, 32'd2990},
{-32'd324, 32'd1211, 32'd8174, -32'd5453},
{-32'd14825, -32'd11342, -32'd14740, -32'd10931},
{-32'd117, 32'd8547, 32'd930, 32'd3477},
{-32'd7204, 32'd3065, -32'd3714, -32'd4972},
{-32'd2028, 32'd6103, -32'd5116, 32'd5619},
{-32'd2562, 32'd3457, -32'd1642, 32'd1381},
{-32'd9066, -32'd7284, 32'd2391, 32'd4707},
{32'd5273, 32'd9083, 32'd4189, -32'd2306},
{-32'd10037, -32'd14287, -32'd6624, -32'd5732},
{-32'd2796, -32'd1478, 32'd4517, -32'd3793},
{-32'd330, -32'd6936, -32'd7289, 32'd1944},
{-32'd2747, -32'd1123, -32'd806, -32'd6124},
{-32'd4295, 32'd7126, -32'd16304, -32'd8548},
{32'd5939, 32'd7936, 32'd4962, 32'd6942},
{32'd11101, 32'd9220, 32'd2019, 32'd12634},
{-32'd6954, -32'd11634, 32'd6584, -32'd7396}
},
{{-32'd1380, 32'd5528, 32'd10934, 32'd3637},
{32'd3067, -32'd1071, -32'd8791, -32'd8542},
{32'd2653, 32'd50, -32'd1873, -32'd4245},
{-32'd5729, -32'd3208, 32'd87, 32'd4646},
{-32'd1290, 32'd105, 32'd10115, 32'd12168},
{32'd9738, 32'd4978, 32'd2849, 32'd7777},
{-32'd2444, -32'd1317, 32'd3056, 32'd8547},
{32'd11860, -32'd2621, -32'd5880, -32'd8972},
{32'd11436, -32'd4253, -32'd2887, -32'd1034},
{-32'd1292, -32'd3510, 32'd4467, 32'd343},
{-32'd1898, -32'd6381, -32'd3199, -32'd4215},
{-32'd10757, -32'd7376, -32'd19151, 32'd1399},
{32'd15027, 32'd18712, -32'd8635, 32'd367},
{32'd5491, -32'd1379, -32'd7456, 32'd8044},
{-32'd4186, 32'd5219, 32'd5229, 32'd2462},
{-32'd5220, 32'd3476, 32'd2862, -32'd2878},
{-32'd5743, 32'd1328, 32'd5450, 32'd3747},
{-32'd7432, 32'd10692, 32'd11869, 32'd7849},
{32'd1626, -32'd21083, 32'd1718, -32'd5923},
{32'd1358, -32'd10045, 32'd6483, -32'd101},
{32'd4603, 32'd1684, 32'd755, 32'd2546},
{32'd6743, -32'd6934, 32'd1803, -32'd11114},
{32'd5602, -32'd1395, -32'd10775, 32'd11712},
{32'd6775, -32'd5240, 32'd144, -32'd1551},
{-32'd11370, 32'd8277, 32'd19477, -32'd479},
{32'd4672, -32'd6197, 32'd968, -32'd4652},
{-32'd5325, -32'd604, 32'd4934, -32'd13643},
{32'd10449, -32'd3066, 32'd17439, 32'd702},
{-32'd4680, 32'd10000, -32'd6656, -32'd3743},
{32'd15908, -32'd754, 32'd2552, -32'd9018},
{32'd7358, 32'd10942, 32'd6296, 32'd10690},
{32'd2577, -32'd9748, 32'd6875, 32'd1977},
{-32'd11173, -32'd4720, 32'd12283, -32'd1678},
{-32'd1443, 32'd6945, 32'd8271, 32'd9769},
{-32'd4015, 32'd3488, 32'd6111, 32'd1209},
{-32'd6048, -32'd1012, 32'd3893, -32'd3261},
{32'd1891, 32'd1960, 32'd1244, 32'd2756},
{-32'd11799, -32'd7766, 32'd8085, 32'd529},
{32'd2692, -32'd1458, 32'd3903, -32'd2194},
{-32'd2265, -32'd2244, -32'd3236, -32'd2560},
{-32'd6330, -32'd814, -32'd18214, -32'd10162},
{-32'd5658, 32'd2108, 32'd5001, -32'd1036},
{-32'd9418, 32'd8338, -32'd15936, 32'd3659},
{32'd518, -32'd4601, -32'd4611, -32'd1449},
{32'd9346, -32'd623, -32'd9983, -32'd238},
{32'd14115, -32'd658, -32'd1439, -32'd1580},
{32'd10418, -32'd969, 32'd2962, 32'd1849},
{-32'd17123, 32'd1287, -32'd3985, 32'd2359},
{32'd2376, 32'd11972, -32'd2186, -32'd2103},
{-32'd5781, -32'd6288, -32'd5246, -32'd833},
{32'd6237, -32'd563, 32'd2695, -32'd12294},
{-32'd8270, -32'd171, 32'd13087, -32'd6347},
{-32'd10682, -32'd10886, -32'd128, -32'd6662},
{-32'd7912, -32'd939, -32'd11638, 32'd16264},
{32'd6292, 32'd15701, 32'd3304, 32'd3085},
{32'd2060, 32'd13763, 32'd5800, -32'd4746},
{32'd16387, -32'd486, 32'd5893, 32'd846},
{-32'd1033, -32'd3802, -32'd2600, -32'd1600},
{32'd1482, -32'd14711, -32'd9400, 32'd829},
{32'd1842, -32'd1013, 32'd2149, -32'd19966},
{32'd3989, -32'd5146, -32'd9371, 32'd1142},
{32'd4641, -32'd5861, 32'd6740, -32'd4598},
{-32'd596, -32'd9196, 32'd129, -32'd1097},
{32'd9894, -32'd2167, -32'd2158, -32'd8166},
{32'd69, -32'd4360, 32'd3573, 32'd5928},
{32'd3766, 32'd8520, 32'd821, 32'd389},
{32'd6514, -32'd8163, -32'd6110, 32'd1781},
{32'd15873, -32'd5748, 32'd1607, 32'd3421},
{-32'd10453, -32'd3502, -32'd5184, -32'd7429},
{32'd4620, 32'd7202, -32'd4360, -32'd12779},
{-32'd241, 32'd849, 32'd6933, -32'd9739},
{-32'd877, 32'd12937, 32'd4177, -32'd486},
{-32'd18005, 32'd4686, 32'd5249, -32'd7705},
{32'd14989, 32'd2559, -32'd7593, -32'd7684},
{32'd6100, 32'd488, -32'd2754, -32'd8946},
{32'd1423, 32'd4312, 32'd6315, 32'd17167},
{-32'd992, 32'd13094, -32'd15413, -32'd1663},
{32'd3021, 32'd2691, -32'd18332, -32'd3939},
{-32'd916, -32'd5003, 32'd95, -32'd2723},
{-32'd9972, -32'd5269, 32'd29923, 32'd5278},
{-32'd3563, -32'd7124, -32'd831, -32'd6040},
{32'd3961, -32'd4501, -32'd6920, -32'd3143},
{-32'd4155, -32'd12823, -32'd3888, -32'd381},
{-32'd5285, 32'd10953, 32'd12041, 32'd16188},
{-32'd8145, -32'd1118, 32'd8130, 32'd11660},
{32'd3777, 32'd3744, -32'd11484, 32'd2864},
{-32'd6790, -32'd7973, 32'd12549, -32'd440},
{-32'd170, -32'd6272, -32'd7754, -32'd1517},
{-32'd3899, -32'd4787, 32'd5681, 32'd3753},
{-32'd5044, 32'd9327, -32'd8497, 32'd3988},
{32'd7363, -32'd2087, 32'd2642, -32'd1021},
{32'd3666, 32'd4833, -32'd5032, 32'd7946},
{-32'd6001, 32'd11400, 32'd5082, -32'd6395},
{32'd3676, 32'd7354, -32'd6180, 32'd1066},
{-32'd6394, 32'd9097, 32'd6157, -32'd3662},
{-32'd4742, -32'd1843, -32'd9140, -32'd2458},
{32'd13844, -32'd515, 32'd4364, -32'd5074},
{32'd1126, 32'd11800, -32'd238, 32'd5462},
{32'd14097, -32'd1498, -32'd2257, 32'd8123},
{-32'd7661, 32'd3632, -32'd3943, -32'd1923},
{-32'd6916, -32'd11655, -32'd954, 32'd11968},
{32'd7406, 32'd18925, 32'd16392, 32'd2684},
{32'd12534, -32'd5645, -32'd925, 32'd16247},
{-32'd5860, 32'd15095, 32'd470, -32'd4963},
{-32'd3720, 32'd2088, -32'd5204, -32'd1491},
{32'd699, 32'd4202, -32'd4581, -32'd6016},
{32'd9973, 32'd6566, -32'd6333, 32'd7331},
{32'd2800, 32'd10874, -32'd1641, 32'd11683},
{32'd3244, -32'd969, -32'd3307, 32'd11227},
{32'd10159, -32'd153, 32'd2913, 32'd722},
{-32'd3109, -32'd557, -32'd1396, 32'd2853},
{-32'd14255, -32'd15718, 32'd272, -32'd12545},
{-32'd1914, 32'd5088, -32'd2028, 32'd9175},
{-32'd24, -32'd9892, -32'd3930, 32'd6061},
{-32'd4529, -32'd159, -32'd4185, 32'd1382},
{32'd3323, -32'd9439, -32'd8882, 32'd12058},
{-32'd14283, -32'd3128, 32'd3433, -32'd8},
{32'd7223, -32'd722, 32'd6426, 32'd1627},
{-32'd4406, 32'd8361, 32'd10321, 32'd4316},
{-32'd444, 32'd1453, -32'd3137, 32'd3886},
{32'd3003, 32'd2109, 32'd1131, 32'd2789},
{-32'd7019, -32'd132, 32'd3498, 32'd5960},
{-32'd962, 32'd15822, -32'd10396, -32'd1273},
{32'd9496, -32'd3653, -32'd7804, 32'd226},
{-32'd13217, -32'd5151, 32'd14605, -32'd3204},
{32'd15109, 32'd4274, 32'd929, -32'd11487},
{-32'd10160, 32'd4415, -32'd2914, -32'd3857},
{32'd2947, -32'd813, 32'd2934, -32'd18276},
{32'd2103, -32'd10229, -32'd7385, -32'd3207},
{-32'd14088, 32'd1090, 32'd11303, -32'd2634},
{32'd4124, 32'd1514, 32'd8638, 32'd825},
{-32'd2057, 32'd2451, -32'd8329, -32'd7483},
{32'd158, 32'd13829, 32'd8598, -32'd2419},
{32'd3154, 32'd3527, -32'd10205, -32'd20210},
{32'd967, -32'd5613, 32'd4521, -32'd7219},
{-32'd4330, 32'd6074, -32'd6206, 32'd289},
{32'd6192, 32'd13174, -32'd5860, 32'd760},
{-32'd1064, 32'd8139, -32'd728, 32'd9107},
{-32'd2246, 32'd6889, 32'd868, 32'd8029},
{-32'd12740, -32'd324, -32'd11665, -32'd8641},
{-32'd12386, -32'd3186, -32'd4178, -32'd13075},
{-32'd123, -32'd4810, -32'd8363, 32'd7187},
{-32'd15892, 32'd8507, 32'd17914, 32'd4643},
{32'd18198, -32'd1272, -32'd13876, 32'd2250},
{-32'd3462, -32'd497, 32'd11073, -32'd4303},
{32'd7874, 32'd8030, 32'd2499, -32'd2851},
{-32'd1580, -32'd11612, 32'd12227, 32'd2091},
{-32'd3938, -32'd3170, -32'd2230, 32'd3650},
{-32'd2145, 32'd6358, 32'd987, -32'd359},
{-32'd9493, 32'd2621, -32'd2612, 32'd2377},
{32'd4470, 32'd1473, 32'd4698, 32'd20929},
{-32'd4051, -32'd2122, -32'd975, -32'd19},
{32'd1117, 32'd11054, 32'd1723, 32'd2095},
{-32'd4213, 32'd1718, 32'd428, -32'd3674},
{32'd9898, -32'd3351, -32'd3098, 32'd5131},
{-32'd3111, -32'd12496, 32'd1813, -32'd415},
{-32'd3041, -32'd5172, -32'd9095, 32'd11356},
{-32'd920, -32'd4195, -32'd2813, -32'd3988},
{32'd6381, -32'd8304, -32'd13962, -32'd3505},
{32'd8504, 32'd3623, -32'd2246, 32'd2062},
{32'd14593, -32'd12453, 32'd3428, -32'd5646},
{-32'd2079, 32'd9024, 32'd2731, -32'd197},
{32'd5620, 32'd2087, -32'd9315, 32'd2581},
{32'd5099, 32'd4817, -32'd6006, 32'd8798},
{-32'd7132, 32'd21034, 32'd2416, -32'd19231},
{32'd2966, -32'd9772, -32'd9535, -32'd3669},
{-32'd518, 32'd8743, 32'd4726, -32'd430},
{32'd3298, -32'd256, -32'd6779, -32'd3421},
{-32'd707, -32'd553, 32'd6449, 32'd14794},
{-32'd14571, -32'd5741, 32'd9915, 32'd15653},
{-32'd3759, 32'd4176, -32'd3047, 32'd8508},
{32'd4552, 32'd4859, 32'd222, 32'd632},
{-32'd459, 32'd58, 32'd2401, 32'd10121},
{-32'd5109, 32'd2026, -32'd371, 32'd9643},
{32'd2695, -32'd6421, -32'd5812, -32'd6162},
{32'd17260, -32'd517, -32'd894, 32'd1405},
{32'd3252, 32'd4805, 32'd12390, 32'd8461},
{32'd14180, -32'd8815, 32'd6344, 32'd7303},
{32'd3850, 32'd9812, 32'd3154, 32'd10870},
{-32'd1172, -32'd9270, -32'd10794, 32'd724},
{-32'd4776, 32'd900, -32'd1672, 32'd5042},
{-32'd4736, -32'd1483, -32'd2281, 32'd7909},
{32'd11019, -32'd9557, -32'd1266, -32'd9107},
{32'd6323, 32'd24092, -32'd2167, -32'd6117},
{32'd10415, 32'd4326, 32'd14472, -32'd1816},
{-32'd12344, 32'd4260, 32'd3229, 32'd3548},
{32'd9409, 32'd6946, 32'd947, -32'd12008},
{32'd514, 32'd15730, 32'd910, 32'd6680},
{32'd11874, -32'd3522, -32'd6246, -32'd253},
{-32'd201, -32'd6985, -32'd17759, 32'd2228},
{-32'd7190, 32'd4054, -32'd4525, 32'd11724},
{32'd1246, 32'd4375, -32'd879, -32'd13567},
{-32'd2087, -32'd10483, -32'd8964, -32'd16239},
{-32'd13359, -32'd410, 32'd4251, -32'd3814},
{32'd5574, -32'd2014, -32'd5309, 32'd11107},
{-32'd17604, -32'd7320, 32'd11593, 32'd4867},
{-32'd20264, -32'd8563, 32'd5689, 32'd18211},
{32'd1297, 32'd5637, 32'd14034, -32'd3201},
{-32'd670, 32'd7563, -32'd11177, -32'd4085},
{32'd7420, 32'd9832, 32'd15454, 32'd468},
{32'd2037, -32'd3731, -32'd6684, 32'd2961},
{-32'd5841, 32'd6274, 32'd2588, -32'd1262},
{32'd12781, -32'd4771, -32'd11848, -32'd9850},
{32'd3303, -32'd1514, -32'd3638, 32'd4956},
{32'd12, 32'd5541, -32'd16197, -32'd10861},
{-32'd3579, -32'd5476, 32'd531, -32'd4507},
{32'd12238, 32'd14295, -32'd3963, -32'd3209},
{-32'd1120, -32'd3126, -32'd2235, -32'd7381},
{32'd8574, 32'd3666, 32'd2996, 32'd5542},
{-32'd161, 32'd5247, 32'd1475, -32'd812},
{-32'd6250, -32'd97, 32'd1123, 32'd7045},
{32'd9105, -32'd563, -32'd2141, 32'd3524},
{-32'd1956, -32'd3792, 32'd12149, 32'd2385},
{-32'd9813, -32'd5502, -32'd4275, -32'd5491},
{32'd5723, -32'd4595, -32'd16637, -32'd291},
{-32'd6627, -32'd11003, -32'd5362, 32'd10442},
{32'd13303, -32'd9244, 32'd6339, 32'd1491},
{-32'd1433, 32'd5785, -32'd6089, -32'd7207},
{32'd17584, -32'd1250, 32'd8635, -32'd993},
{32'd9108, -32'd2699, -32'd2869, -32'd7677},
{32'd14110, 32'd13214, -32'd96, 32'd18399},
{-32'd7172, -32'd9273, -32'd919, -32'd7464},
{32'd16550, 32'd6194, 32'd679, -32'd1648},
{-32'd7105, -32'd12301, 32'd12263, 32'd6988},
{-32'd4047, 32'd3233, -32'd5033, 32'd3715},
{32'd6973, -32'd18435, -32'd10250, 32'd7101},
{-32'd8474, 32'd2947, -32'd16768, 32'd1210},
{32'd1545, -32'd11199, -32'd753, -32'd16684},
{-32'd5767, 32'd9653, 32'd1526, 32'd1378},
{32'd3460, 32'd3291, 32'd7572, -32'd3753},
{-32'd6159, -32'd1006, 32'd924, -32'd8113},
{-32'd13362, 32'd6234, -32'd4405, 32'd3961},
{-32'd2745, -32'd3622, 32'd2252, -32'd1574},
{32'd664, 32'd3481, -32'd2119, 32'd5214},
{32'd11278, 32'd5061, 32'd5098, 32'd9680},
{32'd3309, -32'd19502, 32'd114, 32'd451},
{32'd1153, -32'd4273, -32'd4574, -32'd182},
{32'd5580, -32'd1158, -32'd5688, 32'd741},
{-32'd17596, -32'd2082, 32'd7639, 32'd11546},
{-32'd5288, 32'd5045, -32'd16744, -32'd823},
{-32'd12288, -32'd974, 32'd3383, -32'd1703},
{32'd14227, 32'd5518, -32'd11921, 32'd8260},
{32'd4889, 32'd6849, -32'd3488, -32'd3596},
{32'd6827, 32'd2421, 32'd2499, 32'd10461},
{32'd1734, 32'd1236, -32'd3179, 32'd3674},
{-32'd9160, 32'd2596, 32'd14865, -32'd504},
{-32'd10860, -32'd2532, -32'd1874, 32'd10325},
{-32'd573, -32'd6864, -32'd4311, -32'd18644},
{-32'd4876, -32'd1818, -32'd2077, -32'd6987},
{32'd15271, -32'd8400, 32'd5063, -32'd2502},
{32'd5685, 32'd513, 32'd2961, -32'd5514},
{-32'd20226, 32'd1207, 32'd15887, 32'd7027},
{32'd2257, 32'd4641, 32'd6129, 32'd6240},
{32'd2579, -32'd2614, 32'd5897, -32'd5823},
{32'd11044, -32'd5531, -32'd5528, -32'd993},
{-32'd7249, -32'd8987, -32'd13764, -32'd7485},
{32'd1757, -32'd5730, -32'd7223, -32'd569},
{32'd2886, 32'd15087, -32'd353, -32'd7354},
{-32'd10003, 32'd1855, -32'd1105, -32'd1919},
{32'd13182, -32'd620, 32'd6705, 32'd13668},
{32'd4169, 32'd456, 32'd24058, 32'd6119},
{-32'd2678, -32'd8910, -32'd1833, 32'd12891},
{-32'd10064, 32'd3377, -32'd2134, 32'd5243},
{-32'd8301, 32'd11011, -32'd15617, 32'd4649},
{32'd4368, 32'd271, -32'd821, 32'd6491},
{32'd7343, -32'd7550, -32'd4048, -32'd2278},
{-32'd9662, 32'd4455, 32'd4963, 32'd8215},
{-32'd17445, -32'd811, 32'd7930, 32'd15017},
{-32'd9746, -32'd259, -32'd7640, -32'd2409},
{-32'd189, 32'd758, -32'd799, 32'd5565},
{32'd2394, 32'd406, -32'd2264, 32'd4686},
{32'd4348, 32'd3428, 32'd14467, -32'd1675},
{-32'd4020, -32'd6029, -32'd11505, -32'd15096},
{32'd1251, 32'd5763, 32'd11250, 32'd3927},
{32'd2332, 32'd11551, 32'd6104, -32'd1061},
{32'd1629, -32'd4236, -32'd5223, 32'd4556},
{-32'd2953, 32'd593, 32'd3518, 32'd2155},
{32'd3098, -32'd3101, 32'd10084, 32'd9649},
{32'd2939, 32'd3655, -32'd6425, -32'd751},
{32'd4897, 32'd3905, -32'd3464, 32'd14185},
{-32'd12674, -32'd5204, -32'd666, -32'd5689},
{32'd3938, -32'd2072, -32'd8682, -32'd4176},
{32'd8703, 32'd10104, -32'd7860, 32'd2010},
{32'd525, 32'd62, 32'd7169, -32'd8424},
{-32'd6536, 32'd5320, -32'd10637, -32'd2799},
{-32'd657, -32'd2488, -32'd10897, 32'd112},
{-32'd2594, 32'd3480, -32'd2188, -32'd2946},
{32'd1638, -32'd4547, 32'd3356, 32'd11772},
{32'd2809, -32'd2895, -32'd1535, 32'd18767},
{-32'd18422, -32'd7449, -32'd22833, -32'd5511},
{-32'd4615, 32'd11536, -32'd6534, 32'd5690},
{-32'd6861, 32'd3039, -32'd6911, 32'd1641},
{-32'd239, -32'd942, -32'd8990, -32'd5367},
{32'd7961, -32'd7129, -32'd6787, -32'd7041},
{-32'd5422, -32'd146, -32'd1840, -32'd2773},
{32'd2368, 32'd2554, 32'd523, 32'd21918},
{-32'd15039, 32'd8287, -32'd2643, 32'd3221},
{-32'd549, 32'd4372, 32'd4356, -32'd7386},
{-32'd2924, -32'd402, 32'd14873, -32'd11489},
{-32'd11677, 32'd1004, -32'd568, -32'd5672}
},
{{32'd9666, 32'd3931, 32'd12649, 32'd11684},
{-32'd1202, 32'd2878, -32'd8124, -32'd1},
{32'd9096, -32'd5630, -32'd939, -32'd2935},
{-32'd255, 32'd6777, 32'd3656, -32'd957},
{32'd1114, -32'd1726, 32'd2738, 32'd169},
{-32'd809, 32'd100, -32'd5163, -32'd8435},
{-32'd2455, -32'd6086, 32'd2787, 32'd3025},
{-32'd4232, -32'd5324, 32'd4428, 32'd1478},
{32'd581, -32'd3500, 32'd3361, -32'd716},
{32'd16535, 32'd9923, 32'd4950, 32'd7359},
{32'd868, -32'd3349, -32'd2681, -32'd75},
{-32'd3306, -32'd2484, 32'd7651, -32'd3907},
{-32'd1460, 32'd5578, -32'd3884, 32'd798},
{32'd2216, -32'd2963, -32'd8314, -32'd2687},
{-32'd2333, -32'd8503, 32'd91, -32'd5704},
{-32'd7408, -32'd629, 32'd716, -32'd3589},
{32'd7523, -32'd290, 32'd7404, 32'd1404},
{-32'd823, 32'd6458, 32'd13786, 32'd5947},
{32'd4866, -32'd5221, -32'd7118, -32'd2041},
{32'd4520, 32'd456, 32'd2548, -32'd13194},
{32'd81, 32'd2919, -32'd3089, 32'd4425},
{-32'd9857, 32'd469, -32'd3158, -32'd4967},
{-32'd7907, -32'd1552, -32'd3832, -32'd4376},
{-32'd5543, -32'd6768, -32'd12650, -32'd4700},
{32'd8602, 32'd4703, 32'd798, 32'd8926},
{-32'd2762, 32'd3790, -32'd4314, -32'd6439},
{32'd4447, -32'd28, 32'd9424, 32'd2254},
{-32'd94, -32'd4283, 32'd5207, 32'd1945},
{32'd11750, 32'd13030, 32'd6956, 32'd2180},
{-32'd2226, 32'd240, -32'd7160, -32'd4125},
{32'd1706, -32'd2916, -32'd5277, -32'd1642},
{-32'd16429, -32'd6746, -32'd3190, -32'd467},
{32'd12485, -32'd1063, -32'd2158, 32'd4590},
{-32'd4292, -32'd4973, 32'd2081, 32'd4771},
{32'd8093, 32'd7258, 32'd12547, 32'd5679},
{-32'd1197, -32'd3700, -32'd9317, 32'd2903},
{32'd8268, -32'd2401, 32'd6935, -32'd3650},
{-32'd5578, -32'd2599, 32'd3212, 32'd2403},
{32'd2430, 32'd867, 32'd2280, 32'd3811},
{-32'd894, -32'd975, 32'd2867, -32'd3149},
{32'd5165, -32'd5439, 32'd6710, 32'd267},
{32'd7543, 32'd2210, 32'd1659, 32'd8180},
{32'd1572, -32'd486, 32'd4486, -32'd4141},
{-32'd5420, -32'd8338, -32'd8476, -32'd1459},
{-32'd3561, -32'd718, 32'd10852, -32'd6215},
{-32'd650, -32'd6205, -32'd7249, -32'd2046},
{-32'd7476, -32'd1347, -32'd3929, -32'd2047},
{-32'd6205, 32'd577, -32'd4727, -32'd8105},
{32'd6810, 32'd3643, 32'd957, 32'd8156},
{-32'd2170, -32'd2430, -32'd5068, 32'd3880},
{-32'd3226, 32'd681, 32'd4694, -32'd5883},
{32'd2672, 32'd2844, 32'd3490, 32'd8248},
{-32'd2394, 32'd329, 32'd3321, 32'd52},
{32'd1492, 32'd5280, -32'd14559, 32'd491},
{32'd4533, 32'd4655, 32'd6753, 32'd2829},
{-32'd9746, -32'd2156, -32'd6085, -32'd3130},
{-32'd461, -32'd2511, 32'd11232, 32'd3280},
{-32'd9360, -32'd8701, -32'd9593, -32'd3911},
{-32'd1807, -32'd3640, -32'd6858, -32'd622},
{-32'd3857, -32'd4753, -32'd7156, -32'd9775},
{32'd4845, -32'd2457, -32'd8770, -32'd4493},
{-32'd214, -32'd7256, -32'd2121, 32'd5693},
{-32'd7114, -32'd4642, -32'd7804, -32'd6889},
{32'd584, 32'd32, -32'd690, -32'd2084},
{-32'd3070, 32'd2056, 32'd6000, 32'd1753},
{32'd6989, 32'd6938, 32'd8486, 32'd7726},
{-32'd2318, 32'd1916, 32'd625, -32'd4478},
{-32'd1493, -32'd1001, 32'd2892, -32'd11085},
{32'd4852, 32'd6599, -32'd2806, 32'd2225},
{32'd1772, -32'd959, 32'd1537, -32'd6306},
{-32'd1445, -32'd12512, 32'd2259, -32'd259},
{-32'd2871, -32'd8188, -32'd1018, 32'd6769},
{-32'd1476, -32'd3165, 32'd7452, 32'd249},
{-32'd8203, -32'd4294, -32'd7378, 32'd13703},
{32'd7015, 32'd5638, 32'd5970, -32'd6309},
{32'd8114, -32'd654, -32'd5980, -32'd1544},
{-32'd4362, -32'd7286, -32'd5249, -32'd1416},
{32'd9444, -32'd5803, -32'd12040, 32'd1064},
{32'd784, 32'd5699, -32'd3527, -32'd496},
{32'd8481, 32'd4963, 32'd3295, 32'd3172},
{32'd2720, 32'd7229, 32'd13887, -32'd47},
{32'd2627, 32'd8559, 32'd485, 32'd7495},
{32'd398, -32'd2371, -32'd7378, -32'd7540},
{-32'd4313, 32'd6308, 32'd6174, 32'd471},
{-32'd4201, 32'd2890, -32'd2846, 32'd407},
{-32'd5295, -32'd4570, -32'd4538, -32'd4156},
{32'd2190, 32'd895, 32'd12089, 32'd1902},
{-32'd10173, -32'd3106, -32'd22214, -32'd9044},
{32'd1817, -32'd527, 32'd7428, -32'd11873},
{-32'd8112, -32'd4027, -32'd1098, 32'd1216},
{-32'd876, 32'd190, 32'd3698, 32'd1666},
{-32'd5880, -32'd3087, -32'd8402, 32'd2555},
{32'd6337, 32'd10922, 32'd9734, 32'd8925},
{-32'd1059, 32'd6134, -32'd1647, 32'd6898},
{32'd3844, 32'd2187, 32'd2158, 32'd3643},
{-32'd4823, 32'd3894, 32'd4067, -32'd749},
{32'd8786, 32'd306, 32'd16144, 32'd9527},
{32'd4295, 32'd1599, 32'd2119, 32'd6270},
{-32'd3180, -32'd1578, 32'd470, -32'd5641},
{32'd7671, 32'd9446, 32'd10035, 32'd6881},
{-32'd4027, -32'd2385, 32'd686, 32'd2787},
{-32'd5109, -32'd6292, 32'd3340, 32'd692},
{-32'd898, -32'd2481, 32'd3024, 32'd2967},
{32'd2552, 32'd5221, 32'd1404, -32'd2661},
{-32'd6262, -32'd2608, 32'd2383, 32'd153},
{-32'd1456, -32'd6412, 32'd1273, 32'd2529},
{-32'd1512, -32'd4490, -32'd2647, 32'd2817},
{-32'd2137, -32'd8622, -32'd670, 32'd1772},
{32'd6602, 32'd8096, 32'd8793, 32'd2845},
{-32'd9523, -32'd7350, -32'd2816, -32'd5079},
{32'd6408, -32'd4047, 32'd2493, -32'd3170},
{32'd6466, 32'd6550, 32'd2672, 32'd3523},
{32'd2987, 32'd2397, 32'd5213, -32'd1637},
{-32'd500, -32'd5513, 32'd3973, 32'd8398},
{32'd2253, 32'd842, -32'd5378, -32'd2451},
{32'd2337, 32'd7022, -32'd8266, -32'd325},
{-32'd1414, -32'd2115, 32'd2398, 32'd4134},
{-32'd1498, -32'd290, 32'd6789, 32'd3911},
{32'd1715, -32'd9163, 32'd2992, 32'd8380},
{32'd4286, 32'd5635, -32'd3991, 32'd9411},
{32'd6500, 32'd7058, 32'd5588, 32'd2537},
{32'd12168, 32'd4677, -32'd996, 32'd1176},
{-32'd488, -32'd692, -32'd4680, 32'd7519},
{-32'd2122, -32'd119, -32'd2548, -32'd9829},
{32'd3311, 32'd255, -32'd2751, -32'd1678},
{-32'd6892, -32'd1445, 32'd3254, -32'd3198},
{-32'd933, 32'd1851, -32'd11246, -32'd696},
{-32'd2167, -32'd3750, -32'd4707, -32'd12853},
{-32'd3318, 32'd6587, -32'd1914, -32'd7144},
{32'd6886, 32'd2060, -32'd12291, 32'd1178},
{-32'd1478, -32'd1773, 32'd969, 32'd6348},
{-32'd13615, -32'd1486, 32'd1718, -32'd4156},
{-32'd2604, -32'd662, -32'd3306, -32'd6618},
{-32'd4382, -32'd5524, 32'd5278, -32'd1084},
{32'd4271, -32'd7465, 32'd821, -32'd5211},
{-32'd6186, -32'd1932, 32'd1124, 32'd10547},
{32'd4527, -32'd1335, 32'd3066, 32'd298},
{32'd1137, 32'd5532, 32'd8398, -32'd11187},
{32'd8371, 32'd8907, 32'd11189, 32'd10047},
{32'd6634, -32'd2740, -32'd2636, -32'd930},
{-32'd5090, -32'd8810, -32'd3305, 32'd4121},
{-32'd5457, -32'd1353, 32'd5688, 32'd3039},
{32'd1789, 32'd2019, -32'd349, 32'd3209},
{-32'd3725, -32'd4627, 32'd2444, -32'd6373},
{32'd9960, 32'd1598, -32'd1046, 32'd1456},
{32'd4571, 32'd401, 32'd16553, 32'd6807},
{-32'd4439, -32'd4452, 32'd407, -32'd255},
{-32'd1403, -32'd5095, -32'd165, 32'd3737},
{32'd3156, 32'd6629, -32'd2456, 32'd3137},
{-32'd4391, 32'd5307, -32'd2198, -32'd6025},
{32'd234, -32'd6575, 32'd2260, -32'd6239},
{32'd1260, 32'd4857, 32'd10694, -32'd1386},
{-32'd2133, -32'd3680, 32'd6365, 32'd4483},
{32'd4357, 32'd769, 32'd9001, 32'd255},
{-32'd10205, -32'd9173, -32'd1082, -32'd5057},
{-32'd3661, 32'd2867, -32'd3140, -32'd2876},
{-32'd6293, 32'd7435, 32'd3206, 32'd3025},
{32'd3411, 32'd3659, 32'd7959, 32'd238},
{-32'd2016, 32'd1253, -32'd2061, 32'd1217},
{32'd4749, 32'd6209, -32'd2314, 32'd3437},
{-32'd2103, -32'd1404, 32'd308, -32'd7776},
{32'd2754, 32'd5258, 32'd7918, 32'd3919},
{32'd1796, -32'd900, 32'd652, -32'd325},
{-32'd2827, 32'd4124, 32'd9824, -32'd416},
{-32'd6889, 32'd107, -32'd1221, 32'd2516},
{-32'd8601, 32'd5006, -32'd6445, -32'd6365},
{-32'd3653, 32'd8492, 32'd6618, 32'd1356},
{32'd105, 32'd35, 32'd1104, -32'd7169},
{-32'd2572, -32'd6072, -32'd3532, -32'd6937},
{-32'd8520, -32'd10905, -32'd14659, -32'd7379},
{32'd1530, -32'd3847, 32'd1567, -32'd1370},
{-32'd5795, 32'd5139, -32'd1861, -32'd4226},
{-32'd1154, 32'd5277, 32'd9336, 32'd536},
{-32'd8222, -32'd6139, -32'd2344, 32'd5140},
{-32'd3997, -32'd5621, -32'd9197, 32'd866},
{32'd5951, 32'd5259, -32'd5202, 32'd2005},
{32'd7573, -32'd2322, 32'd690, -32'd4617},
{32'd2931, 32'd5289, 32'd4071, 32'd4582},
{-32'd1926, -32'd3733, 32'd4614, 32'd1674},
{-32'd5598, -32'd6787, 32'd1010, -32'd679},
{-32'd5516, -32'd6644, -32'd4771, 32'd7059},
{-32'd2618, -32'd9894, -32'd1216, 32'd1687},
{-32'd3891, -32'd2695, -32'd9670, -32'd1295},
{32'd6998, -32'd1336, 32'd336, 32'd463},
{-32'd2420, 32'd2001, -32'd903, -32'd3810},
{32'd2163, 32'd3741, 32'd3814, 32'd4250},
{-32'd2192, 32'd1471, 32'd6385, -32'd1045},
{-32'd3663, 32'd5541, 32'd13541, 32'd3886},
{-32'd6310, -32'd614, -32'd3705, -32'd3778},
{-32'd3301, -32'd7978, -32'd12604, -32'd3879},
{-32'd8675, 32'd2943, 32'd5791, 32'd7398},
{-32'd9233, -32'd12416, -32'd14431, -32'd6819},
{-32'd4188, -32'd550, -32'd11158, 32'd455},
{32'd4587, 32'd8079, 32'd7903, 32'd2018},
{32'd3954, 32'd2085, 32'd4089, -32'd158},
{32'd2178, 32'd8754, 32'd5678, 32'd6092},
{-32'd7451, -32'd4232, 32'd5511, 32'd5000},
{32'd2515, 32'd323, -32'd2563, 32'd344},
{32'd2745, 32'd1869, -32'd15489, -32'd13157},
{32'd3124, 32'd2582, 32'd13026, 32'd4036},
{-32'd10925, -32'd6557, -32'd12060, -32'd5653},
{-32'd1106, -32'd205, 32'd7047, 32'd3749},
{-32'd5392, -32'd7261, 32'd1130, -32'd5927},
{-32'd5240, 32'd193, 32'd6965, -32'd2756},
{-32'd3880, 32'd4891, 32'd4112, -32'd4711},
{-32'd248, 32'd8111, 32'd1426, -32'd4319},
{32'd1061, -32'd212, -32'd4164, 32'd3806},
{-32'd6041, -32'd3817, 32'd771, -32'd5397},
{-32'd495, -32'd2150, 32'd8993, -32'd3840},
{32'd7145, 32'd3157, 32'd9561, 32'd4053},
{-32'd2639, 32'd126, -32'd1951, -32'd7196},
{32'd5095, -32'd1837, 32'd7164, 32'd9203},
{32'd1591, -32'd291, 32'd900, -32'd4349},
{32'd13963, 32'd8977, 32'd5675, -32'd397},
{-32'd3435, 32'd6834, 32'd1124, -32'd1160},
{-32'd4168, -32'd4627, -32'd1817, -32'd3613},
{32'd449, -32'd3313, 32'd3040, 32'd5728},
{-32'd805, -32'd1156, -32'd6832, -32'd5675},
{-32'd256, -32'd1436, 32'd12094, 32'd3580},
{-32'd209, -32'd2503, 32'd6677, -32'd1039},
{-32'd7255, -32'd1953, -32'd4115, -32'd5785},
{32'd4172, -32'd3480, -32'd680, 32'd8286},
{32'd5609, -32'd596, 32'd8659, -32'd430},
{32'd2589, -32'd908, 32'd1918, 32'd9685},
{-32'd355, -32'd848, -32'd5580, -32'd267},
{-32'd10713, -32'd468, -32'd6792, -32'd540},
{32'd1553, 32'd4940, -32'd351, 32'd1787},
{32'd2201, 32'd1222, -32'd7711, -32'd5534},
{32'd4127, 32'd7385, 32'd1960, 32'd4283},
{32'd7785, -32'd1184, 32'd8463, 32'd1970},
{-32'd5469, -32'd11142, 32'd1495, -32'd1712},
{-32'd78, -32'd6117, 32'd4922, 32'd2197},
{-32'd2245, 32'd1550, -32'd5889, 32'd6560},
{32'd4578, 32'd116, 32'd4103, 32'd2073},
{32'd2308, 32'd2314, 32'd67, 32'd559},
{32'd1549, -32'd510, -32'd4645, -32'd2393},
{-32'd7487, -32'd1134, 32'd10107, -32'd4201},
{-32'd434, -32'd8089, -32'd3885, -32'd5894},
{-32'd1567, -32'd6494, 32'd553, 32'd4370},
{-32'd917, -32'd4358, -32'd11055, 32'd779},
{32'd695, -32'd3574, -32'd5241, 32'd2116},
{-32'd3370, 32'd10949, -32'd251, 32'd862},
{-32'd7649, -32'd6634, -32'd867, -32'd8514},
{32'd4546, 32'd2629, -32'd5865, -32'd4955},
{32'd10679, 32'd8542, 32'd2961, 32'd10364},
{32'd8239, -32'd3327, 32'd662, -32'd3516},
{-32'd2349, 32'd3165, 32'd5455, -32'd2821},
{-32'd4048, 32'd7306, 32'd187, -32'd2872},
{-32'd4541, -32'd316, 32'd11189, 32'd8279},
{32'd1398, -32'd3081, -32'd328, -32'd274},
{-32'd1245, 32'd3568, -32'd5138, 32'd708},
{32'd2651, 32'd4300, 32'd7602, 32'd6415},
{32'd11461, 32'd3028, 32'd2401, 32'd1077},
{32'd3616, -32'd5844, -32'd1550, -32'd1570},
{-32'd9059, -32'd6184, 32'd1228, -32'd1196},
{32'd573, -32'd4126, 32'd6583, -32'd987},
{32'd1357, 32'd1058, -32'd2640, 32'd2576},
{32'd1243, 32'd1622, 32'd8572, 32'd4498},
{-32'd1523, -32'd2334, -32'd3928, 32'd4869},
{32'd9583, -32'd2435, 32'd8179, 32'd4378},
{32'd7741, 32'd5160, -32'd4564, 32'd408},
{32'd4986, 32'd6198, -32'd6970, 32'd5545},
{32'd3750, 32'd1241, -32'd6164, -32'd6303},
{-32'd6288, 32'd9127, 32'd4187, 32'd1026},
{-32'd8423, -32'd2296, 32'd5594, 32'd5260},
{32'd2272, -32'd2692, -32'd12515, 32'd8001},
{-32'd2592, 32'd5739, -32'd6074, 32'd4263},
{-32'd4703, 32'd2169, 32'd10539, -32'd5728},
{-32'd7443, 32'd1815, -32'd8725, -32'd5325},
{-32'd10430, -32'd3470, 32'd1436, 32'd2545},
{32'd3509, 32'd2694, -32'd4596, -32'd3055},
{32'd3149, 32'd1908, -32'd1648, -32'd264},
{-32'd1738, -32'd8479, -32'd8706, -32'd17},
{-32'd8285, -32'd1102, -32'd7932, -32'd2775},
{-32'd3754, -32'd2334, 32'd5372, 32'd6208},
{32'd1136, -32'd1792, -32'd256, -32'd227},
{32'd13251, 32'd7171, 32'd4852, 32'd9196},
{-32'd5836, 32'd5734, 32'd8307, -32'd1949},
{-32'd4724, -32'd2697, -32'd1929, -32'd7853},
{-32'd3009, -32'd2091, 32'd644, -32'd838},
{32'd7688, 32'd9981, -32'd4547, 32'd2788},
{32'd6138, -32'd4287, 32'd2578, -32'd2961},
{-32'd6544, -32'd2888, 32'd4911, 32'd76},
{-32'd2153, 32'd4472, -32'd8300, -32'd8725},
{32'd11089, 32'd3063, 32'd2095, 32'd2850},
{-32'd4622, -32'd4190, -32'd7991, -32'd11023},
{-32'd4544, 32'd3257, -32'd2969, 32'd835},
{32'd4028, 32'd819, -32'd12310, -32'd1783},
{32'd5726, 32'd2071, 32'd1197, -32'd5004},
{-32'd3192, -32'd5988, -32'd937, 32'd6098},
{32'd2165, -32'd5427, -32'd3702, 32'd590},
{32'd3636, 32'd2294, -32'd5350, 32'd1268},
{-32'd1500, 32'd3642, -32'd3371, -32'd1717},
{32'd2053, 32'd1471, -32'd2830, 32'd820},
{-32'd783, -32'd8006, -32'd4027, -32'd2689},
{32'd3565, 32'd2994, 32'd9483, 32'd2184},
{32'd1528, -32'd825, 32'd2612, 32'd102},
{32'd5683, 32'd13987, 32'd10850, 32'd1565},
{32'd2515, 32'd7687, 32'd4860, -32'd2000},
{-32'd3334, -32'd5853, -32'd10030, -32'd5230}
},
{{32'd3712, 32'd192, 32'd1867, 32'd1046},
{-32'd7670, -32'd3984, 32'd762, 32'd752},
{-32'd438, 32'd912, -32'd4637, -32'd7649},
{32'd11809, 32'd5315, -32'd11559, 32'd948},
{-32'd2889, 32'd674, -32'd3835, -32'd2271},
{32'd8976, -32'd5226, -32'd11499, -32'd7626},
{-32'd984, 32'd1757, -32'd3852, 32'd4349},
{-32'd1761, 32'd1754, 32'd4143, -32'd2729},
{-32'd13920, -32'd3834, -32'd1001, 32'd15650},
{32'd6450, 32'd4932, -32'd7104, 32'd1536},
{32'd3341, -32'd7324, 32'd4761, -32'd12035},
{-32'd4131, -32'd10105, -32'd1464, -32'd19077},
{32'd8350, -32'd1224, 32'd15054, -32'd4558},
{32'd7254, -32'd74, 32'd6653, -32'd7954},
{32'd8294, -32'd6152, -32'd5301, -32'd2281},
{-32'd2318, -32'd17520, 32'd11775, -32'd1327},
{-32'd7938, 32'd671, -32'd542, -32'd6831},
{32'd736, -32'd3319, 32'd4478, -32'd470},
{32'd5709, 32'd4773, 32'd7954, -32'd3928},
{-32'd7616, -32'd3288, -32'd4679, 32'd10051},
{32'd8872, 32'd8413, -32'd7985, -32'd3291},
{32'd2980, 32'd7609, 32'd3528, -32'd7049},
{32'd185, -32'd4394, 32'd4781, 32'd5067},
{32'd6098, -32'd5988, 32'd8260, 32'd11888},
{32'd9518, 32'd3682, -32'd3773, -32'd894},
{32'd10066, 32'd6031, -32'd8591, -32'd918},
{-32'd7230, 32'd10999, -32'd15675, 32'd2273},
{32'd15146, 32'd4215, -32'd4257, 32'd12952},
{-32'd7574, -32'd3715, -32'd1096, 32'd115},
{-32'd5881, -32'd4787, 32'd1773, -32'd1751},
{-32'd4345, -32'd5098, 32'd771, -32'd16639},
{32'd6381, -32'd3266, 32'd6984, 32'd1267},
{-32'd699, 32'd3213, 32'd4973, -32'd2762},
{-32'd3513, -32'd1373, 32'd1485, -32'd9584},
{32'd3811, 32'd2445, -32'd1591, 32'd2947},
{-32'd1413, -32'd5565, 32'd4363, -32'd2067},
{-32'd13032, -32'd8368, 32'd1911, 32'd7452},
{-32'd14978, 32'd647, 32'd7227, 32'd14051},
{32'd5824, -32'd3348, 32'd2671, 32'd3562},
{32'd3312, -32'd2462, 32'd4999, 32'd3504},
{-32'd11214, 32'd411, -32'd2720, 32'd5181},
{-32'd4912, -32'd9859, 32'd9602, 32'd394},
{-32'd1878, -32'd6592, -32'd8171, 32'd4020},
{32'd5533, -32'd6254, 32'd622, 32'd1633},
{-32'd1777, -32'd1697, -32'd3499, -32'd5980},
{32'd2419, -32'd7032, 32'd10966, 32'd3448},
{-32'd2938, -32'd19635, -32'd3493, -32'd3471},
{32'd957, -32'd6328, -32'd5742, -32'd8120},
{32'd2172, 32'd343, 32'd1211, -32'd5583},
{32'd2682, -32'd3438, 32'd7679, 32'd4522},
{-32'd7656, 32'd4045, 32'd1982, -32'd3609},
{32'd7128, -32'd12201, -32'd4784, 32'd5529},
{32'd2473, 32'd8912, 32'd9477, -32'd14893},
{-32'd10803, -32'd6580, 32'd10355, 32'd13432},
{-32'd6401, 32'd5091, -32'd2589, 32'd2481},
{32'd8535, 32'd714, -32'd5801, 32'd2044},
{32'd3973, -32'd84, -32'd1574, 32'd11318},
{32'd3130, -32'd1123, 32'd12165, -32'd402},
{-32'd3486, -32'd4829, 32'd6087, -32'd16450},
{32'd95, 32'd1977, -32'd681, 32'd833},
{-32'd2694, 32'd5584, -32'd6279, -32'd612},
{32'd1130, -32'd2305, 32'd5384, 32'd7130},
{-32'd3039, -32'd8130, 32'd4641, 32'd8697},
{32'd5239, 32'd3771, 32'd2772, 32'd861},
{32'd14122, -32'd1813, -32'd1092, 32'd10949},
{32'd12428, 32'd1705, 32'd626, -32'd3504},
{-32'd1866, 32'd4358, -32'd3975, -32'd6647},
{-32'd1956, -32'd7822, -32'd4225, 32'd4617},
{32'd2160, -32'd8257, -32'd4004, -32'd17469},
{-32'd1942, 32'd4347, 32'd1411, -32'd3132},
{32'd2026, -32'd6942, -32'd906, 32'd8470},
{-32'd4102, -32'd745, -32'd1070, 32'd2557},
{-32'd318, 32'd3801, 32'd4594, -32'd9752},
{32'd43, 32'd7247, 32'd2599, 32'd9568},
{-32'd1745, 32'd12852, 32'd99, -32'd6431},
{-32'd1381, -32'd10445, 32'd6279, 32'd270},
{-32'd5126, -32'd3063, 32'd7471, 32'd13586},
{-32'd10042, -32'd2874, 32'd10404, -32'd12100},
{-32'd6377, -32'd13525, 32'd930, 32'd17988},
{-32'd4883, -32'd1637, -32'd8327, 32'd2670},
{32'd4675, -32'd9468, -32'd6599, 32'd2034},
{32'd3953, 32'd6945, 32'd8352, 32'd935},
{-32'd1414, 32'd2765, 32'd1424, -32'd6096},
{-32'd12473, -32'd4116, -32'd4199, 32'd5623},
{-32'd3147, -32'd4421, 32'd4983, -32'd7865},
{-32'd3993, 32'd1982, -32'd4528, -32'd18587},
{32'd9920, -32'd4071, -32'd3831, 32'd7449},
{-32'd1020, 32'd2565, 32'd5595, 32'd12099},
{-32'd5929, -32'd8018, 32'd5152, -32'd5382},
{-32'd3025, 32'd3931, -32'd12528, -32'd12772},
{32'd11361, 32'd2201, 32'd1553, 32'd9019},
{32'd1468, -32'd1120, 32'd2964, -32'd2726},
{32'd6719, -32'd4510, -32'd2272, -32'd12711},
{-32'd3972, 32'd1101, 32'd5643, 32'd11356},
{32'd6988, 32'd1092, 32'd17809, -32'd165},
{-32'd16646, -32'd4310, -32'd17938, 32'd866},
{32'd10231, 32'd10158, 32'd3511, -32'd3890},
{32'd4404, 32'd2143, 32'd4562, 32'd6383},
{-32'd3032, -32'd1981, 32'd3259, 32'd3214},
{32'd6643, -32'd2681, -32'd2659, -32'd4670},
{32'd2152, -32'd10091, -32'd10146, 32'd13149},
{-32'd20257, 32'd545, -32'd5923, -32'd13876},
{32'd1400, 32'd6821, 32'd1149, 32'd7436},
{-32'd8321, -32'd7088, -32'd11044, 32'd7009},
{32'd3758, 32'd4905, -32'd7347, 32'd2821},
{32'd303, -32'd2584, -32'd3, -32'd4143},
{32'd2414, 32'd10163, -32'd3033, -32'd4141},
{32'd2983, 32'd875, -32'd2939, -32'd2524},
{-32'd5939, 32'd3147, -32'd258, -32'd9114},
{-32'd13542, 32'd609, 32'd1914, 32'd8943},
{-32'd553, -32'd9133, -32'd2721, 32'd4087},
{-32'd2362, 32'd3621, 32'd400, 32'd10045},
{-32'd4026, 32'd29, 32'd10110, -32'd680},
{32'd4881, -32'd138, -32'd1961, 32'd2969},
{-32'd7629, 32'd2982, 32'd8295, -32'd5569},
{-32'd3240, 32'd4977, -32'd8255, 32'd2738},
{32'd458, 32'd395, -32'd2284, -32'd4622},
{32'd6221, 32'd1769, 32'd4909, 32'd8124},
{-32'd12834, 32'd1761, -32'd3963, 32'd13175},
{32'd13080, 32'd2903, 32'd3053, -32'd3825},
{32'd16580, 32'd2653, 32'd2840, -32'd20306},
{32'd2150, 32'd7663, 32'd17780, -32'd8241},
{32'd38, -32'd664, 32'd13095, -32'd4679},
{-32'd687, 32'd5096, 32'd2330, 32'd2623},
{32'd5213, -32'd1164, -32'd5640, -32'd16321},
{32'd4936, -32'd1563, -32'd703, 32'd13822},
{-32'd2908, 32'd11008, -32'd7178, -32'd17744},
{32'd3048, -32'd11920, -32'd1426, -32'd2026},
{-32'd4938, -32'd9407, -32'd2577, 32'd1492},
{32'd1979, -32'd5926, -32'd5500, -32'd588},
{32'd9015, -32'd372, 32'd1011, 32'd2036},
{-32'd17225, -32'd2112, 32'd3254, -32'd748},
{32'd3602, -32'd5020, -32'd13076, 32'd4507},
{-32'd93, -32'd11717, -32'd3637, 32'd11300},
{-32'd7699, -32'd9224, 32'd7421, -32'd4230},
{32'd8419, -32'd8726, 32'd791, -32'd15856},
{-32'd4260, -32'd11125, 32'd1159, 32'd8572},
{-32'd9742, -32'd5558, -32'd3579, 32'd8072},
{32'd5313, 32'd12357, 32'd3116, -32'd3826},
{-32'd12996, -32'd9149, 32'd1432, 32'd6818},
{-32'd1657, 32'd5436, -32'd6993, 32'd14582},
{-32'd4794, 32'd910, -32'd1590, 32'd1755},
{32'd21414, 32'd2308, -32'd5432, -32'd742},
{-32'd9130, -32'd5993, -32'd5782, -32'd5764},
{32'd8702, 32'd2428, -32'd9041, 32'd6448},
{-32'd4186, 32'd650, 32'd1052, 32'd8631},
{32'd7274, -32'd1214, 32'd7121, 32'd149},
{-32'd1125, -32'd589, 32'd2573, -32'd739},
{-32'd4523, 32'd2356, -32'd4870, 32'd5967},
{32'd1829, 32'd15751, -32'd10393, -32'd11435},
{-32'd316, -32'd8480, -32'd1389, -32'd6070},
{-32'd15152, 32'd3601, 32'd601, 32'd11731},
{-32'd8037, 32'd6689, 32'd11432, -32'd6432},
{32'd6206, 32'd5044, -32'd7856, -32'd11753},
{-32'd7054, -32'd9345, 32'd2605, -32'd3234},
{32'd10219, 32'd7830, 32'd3861, -32'd4258},
{-32'd145, -32'd1633, 32'd6692, -32'd6084},
{32'd3430, -32'd8067, -32'd42, -32'd9982},
{32'd5298, -32'd3852, -32'd6252, -32'd676},
{32'd118, -32'd4211, 32'd9165, -32'd5211},
{32'd1178, -32'd3520, 32'd12221, -32'd6367},
{32'd7771, -32'd3985, 32'd6831, -32'd964},
{-32'd4718, -32'd1184, -32'd2517, 32'd6286},
{32'd5795, 32'd5636, 32'd4449, 32'd2966},
{-32'd5931, -32'd8516, -32'd5752, 32'd3174},
{-32'd413, 32'd5359, -32'd8436, 32'd7441},
{32'd2081, -32'd4116, 32'd1799, 32'd1124},
{-32'd5161, -32'd9889, 32'd2969, -32'd7597},
{32'd246, -32'd8088, 32'd12242, 32'd10456},
{32'd11296, -32'd4916, -32'd872, -32'd83},
{32'd1022, -32'd6935, -32'd8688, 32'd2814},
{32'd6097, 32'd2417, -32'd13737, 32'd3686},
{32'd7803, 32'd608, -32'd2662, 32'd6525},
{-32'd2105, -32'd18039, 32'd1153, -32'd728},
{32'd1804, -32'd1106, -32'd2317, -32'd1723},
{32'd7143, 32'd4332, 32'd13562, -32'd9576},
{-32'd793, 32'd4712, -32'd6328, 32'd9756},
{-32'd5408, -32'd1849, 32'd792, -32'd5194},
{32'd4029, 32'd8980, 32'd6355, 32'd7728},
{32'd7904, 32'd3661, -32'd3133, -32'd7844},
{32'd2372, -32'd5565, 32'd4798, 32'd9053},
{-32'd3223, -32'd8329, 32'd3660, -32'd2063},
{-32'd12785, -32'd6554, -32'd818, -32'd5415},
{-32'd4601, -32'd5892, 32'd588, -32'd7228},
{-32'd2051, 32'd1700, -32'd11583, 32'd2232},
{-32'd323, 32'd4484, -32'd7459, -32'd11306},
{32'd4227, -32'd4937, -32'd3832, 32'd10975},
{-32'd4646, 32'd2473, 32'd8840, -32'd11645},
{32'd3571, -32'd551, 32'd5513, 32'd10665},
{32'd9761, -32'd9941, 32'd4815, -32'd3503},
{-32'd7653, 32'd2697, -32'd2902, 32'd11296},
{-32'd8610, -32'd3281, 32'd9077, 32'd6432},
{-32'd9334, -32'd1848, -32'd16325, 32'd5003},
{32'd655, 32'd1638, 32'd2377, 32'd3240},
{-32'd8370, -32'd2242, -32'd1886, -32'd6983},
{32'd1273, -32'd116, -32'd5390, -32'd4456},
{-32'd11539, -32'd345, -32'd15708, 32'd9053},
{-32'd752, -32'd1323, -32'd10923, -32'd2102},
{32'd7194, -32'd9823, -32'd184, -32'd3500},
{-32'd5725, -32'd2974, 32'd943, -32'd2278},
{-32'd6151, -32'd5038, 32'd1890, -32'd731},
{-32'd13407, 32'd6402, -32'd9111, -32'd11835},
{32'd1155, 32'd7089, 32'd2057, 32'd10188},
{32'd7030, 32'd13302, 32'd2566, 32'd7061},
{32'd14313, -32'd15674, -32'd6540, -32'd3525},
{-32'd3133, -32'd7181, 32'd372, 32'd9532},
{-32'd5167, 32'd11838, 32'd3253, 32'd4959},
{32'd3773, -32'd1724, 32'd46, -32'd3879},
{-32'd2081, -32'd6571, 32'd6817, -32'd2599},
{-32'd4047, 32'd3419, 32'd1169, -32'd9038},
{-32'd9489, -32'd9580, 32'd5665, 32'd6411},
{32'd5054, 32'd10101, 32'd859, -32'd2355},
{-32'd11776, -32'd3122, 32'd11318, -32'd2713},
{32'd465, 32'd2421, 32'd4876, -32'd4161},
{32'd11386, 32'd9642, 32'd2969, -32'd887},
{32'd3522, -32'd5441, -32'd473, 32'd4772},
{-32'd6340, 32'd7855, -32'd1339, 32'd18767},
{32'd12746, -32'd5641, -32'd1483, 32'd1940},
{-32'd14016, -32'd561, 32'd4371, 32'd10204},
{32'd4491, 32'd514, -32'd649, 32'd8245},
{32'd1510, -32'd9666, 32'd11650, 32'd12197},
{-32'd16378, 32'd300, -32'd200, 32'd1842},
{-32'd608, 32'd30, 32'd12089, -32'd3415},
{-32'd2361, 32'd14010, 32'd5250, -32'd7251},
{32'd8695, 32'd7799, 32'd8819, -32'd14923},
{32'd3263, 32'd9274, 32'd4623, 32'd7601},
{-32'd7320, -32'd12852, 32'd4562, -32'd11925},
{32'd7267, 32'd3217, -32'd7321, -32'd5519},
{-32'd12955, -32'd4722, -32'd876, 32'd2432},
{32'd14597, 32'd6367, -32'd3435, 32'd15003},
{-32'd3550, -32'd1223, -32'd2109, -32'd4597},
{-32'd9521, -32'd3273, 32'd2411, -32'd3038},
{32'd3919, -32'd2150, 32'd1619, -32'd4574},
{32'd1018, -32'd6080, -32'd10597, -32'd8920},
{32'd13761, -32'd1020, -32'd1408, -32'd5839},
{32'd2354, 32'd5709, -32'd7364, -32'd6720},
{-32'd4506, -32'd822, 32'd4425, -32'd9908},
{32'd8315, 32'd239, -32'd5816, 32'd2005},
{-32'd6133, 32'd99, -32'd6718, -32'd484},
{32'd8172, -32'd9895, -32'd1870, -32'd7141},
{32'd5573, 32'd311, 32'd9806, -32'd4522},
{-32'd1341, 32'd4384, -32'd80, -32'd2974},
{-32'd3110, 32'd170, -32'd8292, 32'd977},
{32'd1473, -32'd1917, 32'd3671, 32'd9560},
{32'd8248, 32'd8144, -32'd1686, -32'd1508},
{-32'd932, -32'd1820, -32'd3805, -32'd3808},
{32'd5123, -32'd4539, 32'd4728, 32'd4255},
{-32'd235, 32'd2679, -32'd8764, -32'd11590},
{32'd2212, 32'd7559, 32'd764, -32'd14882},
{32'd3848, 32'd2157, -32'd5716, 32'd2023},
{-32'd9699, 32'd10793, 32'd13242, 32'd4123},
{32'd8615, -32'd9838, -32'd5659, -32'd7080},
{32'd10525, 32'd830, -32'd1877, -32'd1535},
{32'd4427, 32'd2014, -32'd49, 32'd483},
{-32'd5211, -32'd588, 32'd6313, 32'd9655},
{-32'd2494, -32'd6690, -32'd2988, 32'd11150},
{32'd763, -32'd9069, -32'd16913, 32'd2595},
{32'd8987, 32'd13537, -32'd3180, -32'd12102},
{32'd2371, -32'd1983, -32'd4194, 32'd2911},
{-32'd5956, 32'd5177, 32'd1416, 32'd14097},
{32'd10588, 32'd1799, 32'd1177, 32'd7768},
{32'd14979, -32'd418, 32'd1251, -32'd7147},
{-32'd8116, -32'd14579, -32'd239, -32'd60},
{-32'd4917, -32'd3615, -32'd10242, -32'd13706},
{-32'd6495, 32'd3953, -32'd7045, 32'd15425},
{32'd2059, 32'd2111, 32'd193, 32'd4080},
{32'd16575, 32'd157, 32'd8524, 32'd2998},
{-32'd3920, -32'd1026, 32'd2247, -32'd2913},
{-32'd5206, -32'd13572, -32'd2185, -32'd18679},
{-32'd5069, -32'd9164, -32'd693, 32'd3902},
{-32'd6218, -32'd929, -32'd9746, -32'd7298},
{-32'd16922, -32'd4232, 32'd3969, -32'd6105},
{32'd5654, -32'd3767, -32'd1985, 32'd2797},
{-32'd10357, -32'd3651, 32'd3971, 32'd2057},
{-32'd745, -32'd104, -32'd4472, -32'd13672},
{-32'd2569, -32'd8593, -32'd1243, -32'd1134},
{32'd11673, 32'd8118, -32'd1871, 32'd88},
{32'd382, -32'd4290, 32'd7195, -32'd9535},
{-32'd2758, -32'd7053, 32'd957, -32'd12742},
{32'd4429, 32'd148, 32'd938, -32'd9942},
{32'd7533, 32'd3409, 32'd190, -32'd2652},
{-32'd5219, 32'd5132, 32'd6996, 32'd4988},
{-32'd8287, -32'd212, -32'd4664, -32'd5263},
{32'd18335, -32'd11619, -32'd2028, 32'd15709},
{-32'd1778, -32'd6972, -32'd2140, -32'd6452},
{32'd8988, -32'd2107, 32'd9139, 32'd490},
{32'd558, 32'd13552, 32'd5701, 32'd2453},
{32'd1655, 32'd10742, 32'd9072, 32'd3039},
{32'd9499, -32'd11388, -32'd9514, 32'd20816},
{-32'd51, 32'd3318, 32'd313, -32'd6731},
{-32'd1839, -32'd4311, 32'd16144, -32'd4237},
{32'd10461, 32'd5199, -32'd2568, 32'd2697},
{-32'd7085, 32'd5138, 32'd2175, -32'd8734},
{32'd6474, -32'd1723, 32'd9964, -32'd7330},
{32'd5406, 32'd10449, -32'd2216, -32'd8777},
{-32'd4532, -32'd10660, -32'd5220, -32'd4148},
{32'd3916, -32'd4942, 32'd9551, 32'd597},
{32'd9281, 32'd3640, 32'd4433, -32'd7922},
{-32'd1474, 32'd5168, -32'd9039, 32'd2294},
{32'd7625, -32'd1688, -32'd1649, 32'd6701}
},
{{32'd7928, -32'd8841, 32'd223, -32'd16893},
{-32'd13232, -32'd6882, 32'd1114, 32'd2032},
{-32'd6820, 32'd1500, 32'd8045, 32'd6901},
{32'd7275, -32'd4832, -32'd2437, 32'd10532},
{-32'd3504, 32'd20518, 32'd5698, -32'd1696},
{-32'd6657, 32'd8257, -32'd4791, 32'd3509},
{-32'd4812, 32'd1928, 32'd6633, -32'd1629},
{-32'd1426, -32'd4857, -32'd5935, 32'd9323},
{32'd6042, 32'd13824, 32'd7479, 32'd11041},
{32'd13455, 32'd625, 32'd296, -32'd1914},
{-32'd3469, -32'd263, -32'd1348, 32'd6546},
{32'd1283, -32'd13380, 32'd2326, -32'd12645},
{-32'd7334, -32'd2537, 32'd5496, -32'd1295},
{-32'd197, -32'd966, 32'd3603, -32'd5978},
{32'd1702, -32'd6748, -32'd11317, 32'd1333},
{-32'd4518, -32'd12058, 32'd1000, -32'd12920},
{-32'd205, -32'd4647, -32'd1024, -32'd4664},
{32'd2998, -32'd7105, -32'd4722, 32'd1683},
{32'd7997, -32'd16644, -32'd11578, 32'd18367},
{32'd11866, -32'd5503, 32'd2293, 32'd15968},
{32'd1582, -32'd9384, -32'd7372, 32'd5301},
{-32'd4846, 32'd2721, -32'd9860, 32'd11193},
{-32'd6493, -32'd1395, -32'd10741, 32'd8043},
{-32'd13137, 32'd3251, -32'd7993, 32'd3876},
{32'd7337, -32'd610, -32'd3864, -32'd4973},
{-32'd2616, -32'd7424, 32'd2759, -32'd4979},
{-32'd10193, 32'd4189, 32'd5719, 32'd1328},
{32'd1831, -32'd777, -32'd11627, 32'd6208},
{32'd1885, -32'd17578, 32'd3341, 32'd3742},
{32'd1936, 32'd8781, 32'd10894, -32'd4455},
{32'd1891, -32'd12527, 32'd18, 32'd2476},
{-32'd7537, -32'd6264, 32'd6765, 32'd1086},
{-32'd2715, -32'd2920, 32'd8190, -32'd7327},
{-32'd3439, -32'd12893, 32'd642, -32'd19979},
{32'd4888, 32'd657, -32'd4364, 32'd8545},
{-32'd6477, 32'd8643, 32'd9481, 32'd4394},
{-32'd16239, 32'd3198, 32'd4255, -32'd3126},
{32'd2232, 32'd7094, 32'd6381, -32'd5873},
{32'd1749, -32'd9759, -32'd2971, -32'd11853},
{32'd4955, 32'd2626, -32'd1259, 32'd7775},
{32'd1672, -32'd9217, 32'd4122, 32'd8780},
{32'd12331, 32'd7349, -32'd1289, 32'd4249},
{-32'd13217, -32'd4069, -32'd3708, -32'd8364},
{-32'd4753, -32'd8620, -32'd5697, -32'd11853},
{32'd3108, 32'd1340, 32'd8960, -32'd7110},
{-32'd3697, 32'd1668, 32'd19763, -32'd12552},
{-32'd3017, -32'd7088, 32'd2406, 32'd17169},
{-32'd2472, -32'd16468, 32'd4528, -32'd3007},
{-32'd1335, 32'd4712, -32'd3482, 32'd4106},
{-32'd4997, 32'd6937, -32'd6133, -32'd6176},
{-32'd9464, 32'd5039, 32'd13935, -32'd13757},
{-32'd3230, -32'd1051, -32'd2308, -32'd12395},
{-32'd9866, -32'd16997, -32'd7899, 32'd1552},
{-32'd10080, -32'd7392, -32'd2982, -32'd22097},
{-32'd804, -32'd16039, -32'd7440, 32'd1813},
{32'd7988, 32'd4767, 32'd6351, 32'd10385},
{32'd1421, -32'd7476, -32'd2168, 32'd16550},
{-32'd9361, 32'd2965, -32'd1932, 32'd2023},
{-32'd9222, 32'd370, -32'd659, -32'd4693},
{32'd2183, -32'd3955, 32'd3064, -32'd1527},
{-32'd4482, -32'd5669, 32'd16953, -32'd1404},
{32'd9738, 32'd2828, -32'd1021, 32'd6572},
{-32'd3878, -32'd15, -32'd3992, 32'd7462},
{32'd348, 32'd9767, 32'd18805, 32'd12833},
{32'd6558, -32'd5407, -32'd4867, -32'd11444},
{-32'd182, 32'd6664, -32'd2829, 32'd5723},
{-32'd5596, -32'd6779, 32'd17031, -32'd4126},
{-32'd6959, -32'd4571, -32'd796, -32'd483},
{-32'd8603, -32'd5359, 32'd614, -32'd5865},
{32'd4854, 32'd11653, 32'd2271, 32'd1844},
{-32'd1998, 32'd12953, 32'd1707, -32'd316},
{32'd3773, 32'd539, -32'd1499, -32'd3285},
{-32'd9838, -32'd6144, 32'd2, -32'd4480},
{32'd2289, 32'd3479, 32'd682, 32'd2463},
{32'd153, -32'd8914, 32'd3069, 32'd3404},
{-32'd1340, -32'd5934, -32'd527, -32'd8421},
{-32'd5652, -32'd1778, 32'd7106, -32'd165},
{-32'd10265, -32'd3112, 32'd4726, -32'd6083},
{-32'd3779, 32'd9545, 32'd5160, 32'd2534},
{-32'd4532, -32'd5488, -32'd8432, -32'd10669},
{32'd4005, -32'd1980, 32'd7807, -32'd9449},
{-32'd7620, 32'd5937, 32'd2367, 32'd5739},
{-32'd7709, 32'd5178, 32'd5076, 32'd303},
{32'd6391, -32'd19995, -32'd7079, -32'd5427},
{-32'd7560, -32'd1212, 32'd6231, -32'd13934},
{-32'd5312, -32'd13605, 32'd7927, 32'd2260},
{32'd2482, -32'd10170, -32'd4627, 32'd4614},
{-32'd1450, 32'd7344, -32'd7459, -32'd927},
{32'd12282, -32'd7909, -32'd7467, -32'd10753},
{32'd7658, -32'd8607, -32'd14556, -32'd4026},
{32'd7874, -32'd3765, 32'd6329, -32'd3765},
{-32'd1568, 32'd4596, -32'd3849, 32'd10966},
{32'd2586, 32'd74, -32'd14054, 32'd4761},
{-32'd3168, -32'd11720, 32'd6376, -32'd8237},
{-32'd5279, -32'd5979, -32'd8472, 32'd9776},
{-32'd7879, -32'd4394, 32'd155, 32'd490},
{32'd541, 32'd4457, 32'd4329, 32'd2031},
{-32'd2072, 32'd9609, 32'd7128, -32'd18104},
{-32'd4732, 32'd11980, 32'd4169, 32'd6301},
{32'd10564, 32'd4875, 32'd6168, -32'd3043},
{32'd3744, -32'd12396, -32'd2965, -32'd13731},
{32'd11514, 32'd1861, 32'd115, -32'd4225},
{-32'd6143, -32'd3913, 32'd7625, -32'd3480},
{-32'd10358, -32'd7664, -32'd422, -32'd5314},
{32'd1335, 32'd10793, -32'd11544, -32'd1007},
{32'd423, 32'd10427, 32'd9050, 32'd13043},
{-32'd1483, 32'd2303, 32'd2712, 32'd8657},
{32'd12288, -32'd2614, -32'd8120, -32'd7712},
{32'd2408, 32'd4841, -32'd267, -32'd12159},
{32'd2677, -32'd2940, 32'd3698, -32'd7610},
{32'd444, 32'd12951, -32'd2961, -32'd8626},
{-32'd7565, -32'd2989, -32'd3389, -32'd5359},
{-32'd8172, -32'd6750, -32'd1776, 32'd1080},
{32'd3271, -32'd4027, -32'd6741, -32'd6062},
{-32'd2374, -32'd2010, -32'd2386, 32'd10929},
{-32'd11784, 32'd14257, 32'd3004, 32'd5461},
{32'd13438, -32'd1246, -32'd9698, 32'd11239},
{-32'd4890, -32'd830, 32'd14484, 32'd8024},
{32'd4851, 32'd8138, 32'd10663, 32'd4484},
{-32'd254, -32'd358, -32'd7255, 32'd8177},
{-32'd287, -32'd3779, -32'd6637, -32'd5564},
{-32'd1157, -32'd5817, -32'd17338, -32'd4758},
{-32'd13071, -32'd1193, 32'd1836, -32'd2578},
{-32'd6878, 32'd3450, 32'd1441, 32'd16750},
{-32'd767, 32'd1927, -32'd6867, -32'd5524},
{-32'd6758, -32'd1671, 32'd2813, 32'd3487},
{-32'd2835, 32'd9529, 32'd6250, 32'd6157},
{32'd8569, 32'd7307, 32'd2161, 32'd2798},
{32'd996, -32'd4410, -32'd2965, 32'd4764},
{32'd4462, -32'd6923, -32'd402, -32'd19625},
{-32'd5807, 32'd8968, 32'd5425, 32'd13927},
{-32'd10644, 32'd6389, 32'd4380, -32'd11743},
{-32'd7541, -32'd5794, 32'd1140, -32'd4008},
{-32'd11443, 32'd16970, 32'd10806, -32'd529},
{32'd1631, 32'd14751, -32'd5389, 32'd25552},
{32'd242, 32'd6212, -32'd1027, -32'd6044},
{32'd2022, -32'd5487, 32'd9380, 32'd6655},
{32'd8780, 32'd12393, 32'd9893, -32'd2227},
{32'd4137, -32'd2469, 32'd6123, 32'd600},
{-32'd11459, 32'd819, 32'd4398, 32'd4483},
{-32'd6493, 32'd10219, 32'd4144, -32'd3445},
{32'd2134, -32'd1301, 32'd14611, -32'd2966},
{32'd5495, -32'd14367, -32'd12111, 32'd3403},
{-32'd3518, -32'd10252, 32'd4290, -32'd6891},
{32'd21, -32'd17180, -32'd7168, -32'd1521},
{-32'd8637, 32'd10327, 32'd6893, -32'd5571},
{-32'd2107, 32'd3509, 32'd2327, 32'd1633},
{32'd5619, 32'd7510, 32'd3259, -32'd4379},
{32'd3693, 32'd12094, 32'd6100, 32'd14731},
{-32'd3387, -32'd10013, -32'd7621, -32'd2844},
{-32'd9814, -32'd12678, -32'd11116, -32'd9080},
{32'd11553, 32'd4153, 32'd10777, -32'd4974},
{-32'd647, 32'd12526, -32'd3023, -32'd10616},
{-32'd4970, -32'd4844, 32'd7004, 32'd3593},
{-32'd10135, 32'd17248, -32'd809, 32'd12917},
{-32'd2967, 32'd5813, 32'd2214, 32'd1246},
{32'd15088, 32'd3246, -32'd7751, 32'd9676},
{32'd16326, -32'd14714, -32'd8474, 32'd6919},
{-32'd14022, -32'd16117, 32'd315, -32'd13001},
{32'd4352, 32'd2086, 32'd1273, -32'd5523},
{32'd7767, -32'd1092, 32'd6306, -32'd11737},
{32'd3154, -32'd5149, 32'd1115, -32'd7592},
{-32'd14427, -32'd7384, -32'd221, -32'd1973},
{32'd3876, 32'd5912, -32'd5242, -32'd5443},
{-32'd3604, 32'd8150, -32'd5432, -32'd4341},
{32'd990, 32'd3577, 32'd5655, -32'd10355},
{-32'd5717, -32'd6718, 32'd300, -32'd6434},
{-32'd387, -32'd9333, 32'd3491, 32'd3194},
{-32'd13301, -32'd2071, 32'd4000, 32'd2513},
{32'd148, -32'd12436, -32'd14910, 32'd934},
{32'd7065, -32'd37, -32'd1588, -32'd3067},
{32'd2997, 32'd6800, -32'd9445, 32'd7749},
{32'd7994, 32'd3224, -32'd2204, 32'd3280},
{-32'd15967, -32'd9386, -32'd5275, 32'd14281},
{32'd7305, 32'd2737, -32'd2012, 32'd13037},
{32'd4224, 32'd656, 32'd7565, -32'd10374},
{-32'd5018, 32'd8016, -32'd4584, -32'd10432},
{32'd7899, -32'd1008, 32'd3586, -32'd4802},
{-32'd4491, 32'd19298, 32'd3678, 32'd2447},
{-32'd3382, -32'd8645, -32'd477, -32'd8652},
{32'd2415, -32'd8491, 32'd5480, -32'd15912},
{-32'd5819, -32'd7407, 32'd672, -32'd15117},
{32'd4749, -32'd14780, 32'd2342, 32'd3989},
{32'd670, -32'd2750, -32'd7597, -32'd10338},
{32'd1022, 32'd7335, -32'd13927, 32'd13141},
{32'd8927, 32'd3010, -32'd5980, 32'd5073},
{32'd11191, 32'd15104, 32'd11065, 32'd17665},
{32'd2615, 32'd6289, 32'd19114, -32'd14353},
{32'd5434, 32'd16568, 32'd7129, 32'd1586},
{32'd3690, -32'd8968, 32'd7577, -32'd1801},
{-32'd3962, 32'd4642, -32'd3667, 32'd539},
{-32'd7843, 32'd6164, 32'd11405, -32'd126},
{-32'd5142, -32'd2836, -32'd10795, 32'd4448},
{-32'd1166, 32'd7032, -32'd1476, 32'd5100},
{32'd11881, -32'd157, 32'd1394, -32'd11509},
{32'd6484, -32'd2420, -32'd11412, -32'd9606},
{32'd1663, -32'd2043, -32'd13427, 32'd9058},
{-32'd6600, -32'd947, 32'd5273, -32'd6713},
{32'd8107, 32'd4214, 32'd9894, 32'd2108},
{-32'd8092, -32'd382, 32'd763, -32'd13438},
{-32'd3372, 32'd2940, -32'd2966, 32'd5340},
{-32'd5153, 32'd172, -32'd1042, 32'd989},
{32'd2798, 32'd24717, 32'd16639, -32'd3619},
{32'd436, 32'd10665, 32'd8089, 32'd6608},
{-32'd6023, -32'd20063, 32'd3989, -32'd5975},
{-32'd1134, -32'd13354, 32'd8596, 32'd1309},
{32'd13270, 32'd16931, -32'd868, 32'd4682},
{32'd596, -32'd8573, -32'd374, -32'd7540},
{32'd7350, -32'd4004, -32'd9715, -32'd6002},
{32'd3950, -32'd5517, -32'd4217, -32'd14359},
{-32'd6581, -32'd14058, 32'd6515, -32'd7602},
{32'd12560, -32'd7989, 32'd2540, -32'd21252},
{32'd4288, 32'd4106, 32'd5115, 32'd2876},
{32'd6972, 32'd3423, 32'd5347, -32'd2609},
{-32'd9542, -32'd13386, -32'd1639, 32'd5125},
{-32'd665, -32'd4519, -32'd829, 32'd5893},
{32'd660, 32'd12909, 32'd11229, 32'd8530},
{-32'd5098, -32'd8986, -32'd2558, 32'd3506},
{-32'd1860, 32'd3913, 32'd15693, 32'd61},
{-32'd7432, 32'd2890, 32'd4968, 32'd180},
{32'd6242, 32'd7019, 32'd9028, -32'd7096},
{-32'd166, 32'd15593, -32'd3470, -32'd2892},
{-32'd95, 32'd15947, -32'd7102, -32'd749},
{-32'd2136, -32'd7250, 32'd2001, -32'd2170},
{32'd2873, -32'd5028, -32'd7087, -32'd1635},
{-32'd4162, -32'd9299, -32'd1386, 32'd3806},
{32'd4007, -32'd12225, 32'd9290, 32'd4934},
{-32'd2156, -32'd7214, -32'd872, 32'd1438},
{32'd1569, -32'd7781, 32'd3380, 32'd3547},
{32'd4112, -32'd999, 32'd2055, -32'd2240},
{-32'd1415, 32'd9003, -32'd5431, 32'd8086},
{-32'd5937, -32'd3820, 32'd5795, -32'd3167},
{-32'd713, -32'd2233, -32'd3862, 32'd2696},
{32'd9955, -32'd5452, 32'd325, -32'd10012},
{32'd1201, -32'd4974, 32'd7188, -32'd4164},
{-32'd8273, 32'd993, 32'd8957, 32'd4571},
{-32'd1695, 32'd9896, 32'd3276, -32'd6447},
{-32'd17442, 32'd5746, 32'd2561, 32'd14734},
{32'd6805, 32'd9835, -32'd12044, -32'd1332},
{-32'd1524, 32'd334, -32'd3451, 32'd13325},
{32'd3860, -32'd852, 32'd5540, 32'd10807},
{32'd13521, -32'd6006, 32'd844, 32'd2974},
{-32'd9210, -32'd15214, -32'd7446, 32'd9877},
{32'd8245, 32'd4531, -32'd480, -32'd5636},
{32'd3614, 32'd1785, -32'd4145, -32'd538},
{-32'd5195, -32'd969, -32'd4812, 32'd10282},
{-32'd8194, -32'd6760, 32'd8214, -32'd6143},
{32'd5540, 32'd3502, -32'd3820, 32'd11160},
{32'd5816, -32'd18416, -32'd6750, 32'd6412},
{-32'd234, 32'd40, 32'd18, 32'd2277},
{32'd6399, 32'd7009, 32'd6969, -32'd9195},
{32'd7749, -32'd8375, -32'd9757, 32'd16671},
{32'd92, 32'd7689, 32'd4908, -32'd21213},
{-32'd8506, 32'd1718, -32'd4752, 32'd9327},
{-32'd6406, 32'd3187, 32'd12580, -32'd3264},
{-32'd3297, -32'd5872, 32'd7117, 32'd13569},
{32'd2649, 32'd5444, -32'd335, -32'd2009},
{32'd6346, 32'd11375, -32'd5950, -32'd515},
{-32'd7831, -32'd5818, -32'd7667, 32'd16},
{32'd767, 32'd5295, 32'd8459, -32'd20161},
{32'd9211, 32'd939, -32'd3069, 32'd11581},
{32'd685, -32'd7845, -32'd11654, -32'd15400},
{-32'd9741, -32'd20770, -32'd5719, 32'd986},
{-32'd7193, -32'd11725, -32'd6734, -32'd1751},
{32'd1234, 32'd7754, 32'd2356, -32'd10141},
{32'd11384, 32'd1558, 32'd6866, -32'd5852},
{32'd134, 32'd10486, -32'd8674, 32'd13122},
{-32'd859, 32'd4187, -32'd18164, -32'd5182},
{32'd4538, -32'd2632, -32'd10605, 32'd7095},
{-32'd775, -32'd13085, 32'd995, 32'd499},
{-32'd5963, -32'd9944, 32'd284, -32'd6683},
{-32'd2244, 32'd6299, -32'd10578, 32'd1232},
{-32'd5989, -32'd463, 32'd7569, -32'd3952},
{32'd2587, 32'd12420, 32'd14540, -32'd3243},
{32'd5666, 32'd4646, 32'd2009, 32'd8312},
{-32'd10088, -32'd4777, -32'd716, -32'd7437},
{32'd10179, -32'd896, 32'd23, -32'd2739},
{-32'd3297, 32'd9147, -32'd654, 32'd2949},
{-32'd4225, -32'd8672, -32'd8203, -32'd4742},
{-32'd1783, -32'd25165, -32'd5150, -32'd7612},
{32'd7449, 32'd26, -32'd1619, -32'd4044},
{32'd4803, 32'd23216, -32'd3118, 32'd9796},
{32'd518, 32'd12817, 32'd7054, 32'd1963},
{-32'd2834, 32'd3632, 32'd4821, 32'd18823},
{-32'd861, -32'd11379, -32'd8456, -32'd14918},
{-32'd2176, -32'd9934, 32'd850, -32'd4017},
{32'd3575, 32'd2298, -32'd5006, -32'd5363},
{-32'd5158, -32'd8689, -32'd8460, -32'd10111},
{32'd12091, -32'd12537, -32'd75, 32'd1629},
{-32'd3158, -32'd11891, -32'd7685, 32'd3658},
{-32'd7484, 32'd7994, 32'd8596, 32'd3661},
{32'd6288, 32'd11958, -32'd9189, 32'd1509},
{32'd7246, -32'd7165, -32'd352, -32'd6732},
{32'd14187, -32'd4207, 32'd8886, -32'd13828},
{32'd7350, 32'd25, -32'd5110, 32'd5156},
{-32'd4696, -32'd9170, -32'd4398, -32'd17021},
{-32'd5942, -32'd14678, -32'd2711, -32'd2164},
{32'd12504, 32'd3835, -32'd3408, 32'd8978},
{32'd7411, -32'd5502, -32'd7591, 32'd1493},
{-32'd3028, -32'd4070, -32'd5442, -32'd5729}
},
{{32'd3964, 32'd500, 32'd3852, -32'd8608},
{32'd24, -32'd5217, -32'd756, -32'd2889},
{32'd7535, -32'd557, 32'd266, 32'd2096},
{-32'd1212, -32'd2686, 32'd2984, -32'd3615},
{32'd1170, -32'd8381, 32'd4558, 32'd824},
{-32'd1262, 32'd3981, -32'd10700, -32'd499},
{32'd12893, -32'd74, 32'd6744, 32'd3287},
{32'd78, -32'd10766, -32'd3009, -32'd4641},
{-32'd5980, 32'd2379, -32'd2256, 32'd850},
{32'd11055, 32'd9491, 32'd9913, 32'd4270},
{-32'd5415, 32'd805, -32'd2088, 32'd7268},
{32'd12278, 32'd5519, -32'd5781, -32'd8257},
{-32'd5928, 32'd1736, -32'd6909, 32'd4344},
{32'd828, -32'd8115, -32'd297, -32'd6600},
{-32'd3977, -32'd8952, 32'd473, -32'd8793},
{-32'd7462, 32'd120, -32'd4308, -32'd2583},
{32'd1552, -32'd399, 32'd2659, -32'd7167},
{32'd1801, -32'd7378, 32'd734, -32'd4173},
{32'd2174, -32'd3629, 32'd4057, -32'd3158},
{32'd7892, -32'd3140, 32'd9380, -32'd2185},
{32'd2110, -32'd4676, 32'd10844, -32'd3851},
{-32'd1807, -32'd1506, -32'd1409, -32'd2954},
{-32'd3594, -32'd8360, 32'd1582, -32'd8455},
{-32'd3584, 32'd952, -32'd14011, 32'd216},
{32'd4477, 32'd3211, 32'd1898, -32'd2181},
{32'd9417, -32'd7042, 32'd6049, 32'd6249},
{-32'd638, 32'd5793, -32'd7774, 32'd10606},
{32'd7123, 32'd1337, 32'd1832, 32'd12475},
{-32'd1793, 32'd8996, -32'd958, 32'd4298},
{32'd5245, -32'd5352, -32'd3119, -32'd9554},
{-32'd5623, -32'd4976, -32'd404, -32'd10294},
{-32'd4119, -32'd12708, -32'd3308, 32'd4279},
{-32'd5883, 32'd3370, 32'd2599, -32'd700},
{32'd4469, -32'd5504, -32'd6496, -32'd432},
{32'd7364, 32'd2346, 32'd7444, 32'd2965},
{-32'd182, 32'd2559, -32'd8819, 32'd734},
{32'd7109, -32'd4486, -32'd1810, 32'd12849},
{-32'd2843, 32'd4680, 32'd2313, -32'd5085},
{32'd9980, -32'd1776, -32'd2429, 32'd361},
{32'd5558, 32'd11232, 32'd3860, 32'd4361},
{32'd812, 32'd5521, 32'd1986, -32'd3852},
{32'd2420, -32'd3070, 32'd3437, 32'd6791},
{32'd8225, 32'd4365, 32'd3135, -32'd3224},
{-32'd4114, -32'd261, -32'd834, -32'd5735},
{-32'd3739, 32'd162, -32'd2505, 32'd6358},
{32'd3435, 32'd10836, 32'd3900, 32'd3112},
{-32'd10232, -32'd6009, -32'd10163, 32'd2791},
{32'd10673, 32'd365, -32'd10979, -32'd5385},
{32'd9887, 32'd2738, 32'd6506, 32'd2623},
{32'd10077, -32'd7585, 32'd21403, -32'd1383},
{-32'd3380, 32'd6907, -32'd1031, 32'd4794},
{32'd10727, -32'd1555, -32'd5957, -32'd7349},
{-32'd3144, -32'd7343, 32'd1219, 32'd1006},
{-32'd2498, -32'd6433, 32'd7694, -32'd13235},
{-32'd8812, 32'd7040, -32'd4045, -32'd379},
{-32'd5496, -32'd3873, -32'd3574, -32'd2120},
{-32'd719, -32'd1674, 32'd8529, -32'd2724},
{-32'd3120, -32'd4772, -32'd5473, 32'd85},
{-32'd4395, 32'd612, 32'd2381, -32'd13935},
{32'd5673, 32'd5065, 32'd1126, -32'd6568},
{-32'd3043, -32'd1595, 32'd2985, -32'd1438},
{-32'd5416, -32'd3475, -32'd286, 32'd1462},
{-32'd11388, -32'd2535, -32'd8279, 32'd1786},
{32'd723, -32'd6922, 32'd2183, -32'd574},
{32'd4356, -32'd638, 32'd4111, -32'd2572},
{32'd5592, -32'd2632, 32'd3725, 32'd5576},
{32'd7602, 32'd6064, 32'd1678, 32'd1629},
{-32'd5733, -32'd9585, 32'd4142, 32'd578},
{32'd1521, -32'd185, -32'd1664, -32'd3721},
{-32'd749, 32'd2154, 32'd432, -32'd1609},
{-32'd4187, 32'd1392, -32'd10441, -32'd6675},
{-32'd4808, -32'd3462, -32'd8554, 32'd5031},
{32'd1357, 32'd1378, -32'd1624, -32'd5310},
{32'd8917, 32'd2390, 32'd4092, -32'd4612},
{-32'd1129, 32'd2796, 32'd1269, 32'd2161},
{32'd2315, 32'd4808, 32'd931, -32'd13832},
{32'd2160, -32'd142, 32'd2097, -32'd6114},
{-32'd8885, -32'd4543, -32'd2605, -32'd1176},
{32'd7965, 32'd4905, -32'd1275, 32'd5049},
{-32'd3511, 32'd4334, -32'd4017, 32'd4708},
{32'd5194, -32'd3749, 32'd9019, 32'd9709},
{32'd9508, 32'd4541, 32'd4499, 32'd1532},
{32'd1856, -32'd1960, -32'd1321, -32'd5435},
{-32'd1434, -32'd410, 32'd1747, -32'd6969},
{-32'd8077, 32'd2688, -32'd9804, -32'd8367},
{-32'd1143, -32'd840, 32'd8711, 32'd3149},
{32'd11184, 32'd4096, 32'd3821, 32'd1295},
{-32'd14319, -32'd4688, -32'd3477, 32'd1267},
{-32'd3523, -32'd503, -32'd4402, -32'd744},
{-32'd8918, -32'd461, -32'd7179, -32'd7762},
{32'd7105, 32'd4160, 32'd9096, 32'd4286},
{-32'd1025, -32'd11421, 32'd3796, -32'd407},
{32'd535, 32'd5574, 32'd1771, 32'd2875},
{32'd2893, 32'd1115, -32'd767, 32'd3836},
{-32'd8250, -32'd4531, 32'd70, -32'd286},
{-32'd14722, -32'd9870, 32'd6669, -32'd3105},
{-32'd626, 32'd703, 32'd4938, 32'd3676},
{-32'd4116, 32'd10854, -32'd7588, -32'd5658},
{-32'd5785, -32'd8278, 32'd5339, 32'd4250},
{32'd14339, 32'd9742, 32'd3467, 32'd3064},
{32'd895, 32'd1844, 32'd797, 32'd10698},
{32'd3372, -32'd229, 32'd3350, -32'd1812},
{32'd1348, -32'd915, 32'd645, -32'd1930},
{32'd2883, 32'd7924, 32'd1922, -32'd3997},
{-32'd10520, 32'd2508, 32'd2436, -32'd7281},
{32'd4280, -32'd2870, 32'd3796, -32'd3896},
{-32'd4934, 32'd2725, 32'd1071, 32'd3948},
{-32'd3855, -32'd277, 32'd85, -32'd8490},
{-32'd3848, 32'd8497, 32'd1052, 32'd7996},
{-32'd11061, 32'd1720, -32'd2797, -32'd4267},
{32'd2018, -32'd2794, -32'd1715, -32'd804},
{32'd7068, 32'd4168, -32'd1181, 32'd2327},
{-32'd4178, -32'd858, 32'd7309, -32'd2981},
{32'd4088, -32'd365, 32'd2431, 32'd3971},
{32'd1368, 32'd6838, -32'd5808, -32'd10639},
{-32'd5473, -32'd3373, 32'd198, -32'd3437},
{32'd6564, 32'd4371, 32'd2484, -32'd3451},
{32'd5248, -32'd3018, -32'd2943, 32'd1037},
{32'd5974, -32'd578, -32'd1962, -32'd2392},
{32'd4957, 32'd3312, 32'd2379, -32'd4142},
{32'd7366, 32'd1985, -32'd868, -32'd6566},
{32'd1924, 32'd1448, -32'd77, -32'd985},
{32'd12706, 32'd6367, 32'd2675, -32'd2275},
{-32'd4184, -32'd6448, -32'd1169, -32'd4737},
{-32'd3536, -32'd1516, -32'd7852, -32'd6431},
{-32'd7127, 32'd6223, 32'd5222, 32'd5746},
{-32'd12096, 32'd9440, -32'd9826, -32'd6428},
{32'd7116, -32'd5896, 32'd2531, -32'd7474},
{-32'd2017, 32'd6526, -32'd4163, 32'd1591},
{-32'd13336, -32'd3124, -32'd1207, -32'd4706},
{-32'd6662, 32'd1205, -32'd3769, -32'd5880},
{-32'd3524, 32'd232, -32'd6966, 32'd3037},
{-32'd5370, -32'd602, -32'd799, -32'd3937},
{32'd9662, -32'd3201, -32'd5170, 32'd12666},
{32'd7022, -32'd4547, -32'd67, -32'd2769},
{-32'd7188, 32'd2682, -32'd669, -32'd7033},
{-32'd7225, 32'd912, -32'd2432, -32'd2533},
{-32'd1534, 32'd2156, 32'd2461, 32'd6350},
{-32'd8197, -32'd6133, 32'd9390, -32'd4935},
{-32'd4196, 32'd1248, -32'd275, 32'd6944},
{-32'd4890, 32'd1959, -32'd3080, 32'd2979},
{-32'd2444, -32'd5273, -32'd8986, 32'd1120},
{32'd7295, -32'd3760, -32'd859, -32'd3595},
{32'd22, -32'd3830, 32'd11000, 32'd8000},
{32'd8202, 32'd7636, 32'd2314, -32'd3515},
{32'd6195, -32'd5674, 32'd4129, 32'd7995},
{-32'd6628, -32'd1315, 32'd2189, -32'd1870},
{32'd3406, -32'd914, 32'd4694, -32'd6945},
{32'd2384, 32'd1551, 32'd1228, -32'd2840},
{32'd1730, -32'd2800, -32'd3888, -32'd6107},
{-32'd2978, -32'd5077, -32'd3474, -32'd3854},
{-32'd3507, 32'd3964, 32'd782, -32'd7864},
{-32'd7153, 32'd1397, -32'd2481, 32'd331},
{-32'd5266, 32'd4396, 32'd1319, 32'd3595},
{-32'd9538, -32'd1580, -32'd6885, 32'd1446},
{32'd4442, -32'd7060, 32'd6865, 32'd899},
{32'd2280, 32'd4940, 32'd9379, -32'd5724},
{32'd3246, -32'd3718, 32'd11613, -32'd3528},
{-32'd9040, -32'd4499, 32'd14343, -32'd6731},
{32'd8129, -32'd695, -32'd116, 32'd227},
{32'd1942, -32'd7869, 32'd34, 32'd3163},
{32'd3433, 32'd2498, -32'd3003, -32'd3994},
{-32'd771, -32'd5652, -32'd9520, 32'd1123},
{32'd10002, 32'd1601, 32'd7908, -32'd1269},
{-32'd271, 32'd15583, -32'd8193, 32'd6634},
{-32'd11699, -32'd9342, 32'd1544, -32'd4180},
{-32'd4008, 32'd3625, 32'd2165, 32'd3923},
{-32'd4227, 32'd5770, -32'd6912, -32'd6362},
{-32'd34, 32'd4885, -32'd803, 32'd1159},
{-32'd6037, -32'd2834, -32'd9562, -32'd3429},
{-32'd3780, 32'd1574, -32'd9919, -32'd2104},
{-32'd97, -32'd2408, -32'd2214, 32'd5176},
{32'd7439, 32'd3233, 32'd8307, 32'd3393},
{-32'd4646, -32'd9608, -32'd581, 32'd2687},
{-32'd1043, -32'd4231, -32'd1538, -32'd4596},
{-32'd4139, 32'd2680, 32'd758, -32'd6443},
{-32'd2752, 32'd4256, 32'd2435, 32'd1780},
{32'd213, 32'd1399, -32'd1410, -32'd8122},
{32'd9579, 32'd5506, -32'd3817, -32'd13965},
{-32'd396, 32'd1322, -32'd8550, -32'd1671},
{32'd2832, -32'd244, -32'd5327, -32'd11919},
{-32'd6357, -32'd2877, -32'd476, -32'd2407},
{32'd1709, -32'd8350, -32'd1962, -32'd782},
{-32'd5741, -32'd171, -32'd9849, -32'd1126},
{-32'd8476, 32'd4615, -32'd1323, -32'd1496},
{-32'd2236, -32'd10648, 32'd1374, -32'd5422},
{32'd6827, -32'd2562, 32'd2897, 32'd1855},
{32'd9911, 32'd6988, 32'd1088, -32'd7238},
{-32'd12013, -32'd4830, -32'd2403, 32'd1353},
{-32'd2157, 32'd546, 32'd12, -32'd3948},
{32'd4502, -32'd4561, -32'd1133, -32'd3307},
{-32'd8297, -32'd2501, -32'd19450, -32'd1232},
{32'd2111, 32'd4127, -32'd6834, -32'd158},
{32'd3792, -32'd596, 32'd4399, 32'd7585},
{32'd8786, -32'd976, -32'd4201, -32'd2594},
{32'd4230, 32'd2478, 32'd6056, 32'd7973},
{32'd9885, -32'd10535, -32'd250, -32'd2123},
{32'd4062, 32'd4946, 32'd1226, 32'd1107},
{-32'd788, -32'd7605, -32'd2228, -32'd4644},
{-32'd3630, 32'd433, 32'd3959, 32'd4861},
{-32'd6125, -32'd1568, -32'd4974, -32'd2007},
{-32'd6467, 32'd2049, -32'd5769, 32'd6197},
{-32'd5168, 32'd410, -32'd2784, 32'd7466},
{-32'd564, 32'd3445, 32'd3610, 32'd13322},
{32'd412, -32'd887, -32'd4064, -32'd4253},
{32'd1730, 32'd5814, 32'd2865, -32'd2037},
{32'd3989, 32'd2059, 32'd5686, 32'd1675},
{-32'd4544, 32'd3110, -32'd8073, -32'd7483},
{32'd3273, -32'd1202, -32'd122, 32'd5937},
{32'd7209, 32'd7518, -32'd4006, 32'd2360},
{-32'd1724, -32'd1874, -32'd1601, -32'd5},
{32'd3530, -32'd3028, 32'd9374, -32'd4537},
{-32'd2290, -32'd2287, -32'd3465, -32'd4417},
{-32'd45, -32'd2757, -32'd619, 32'd4071},
{-32'd7366, -32'd2557, 32'd1651, 32'd5642},
{-32'd3060, 32'd627, -32'd2372, -32'd1955},
{-32'd684, -32'd2109, 32'd6902, 32'd8090},
{32'd5075, 32'd101, -32'd7664, -32'd5764},
{32'd1151, 32'd7450, -32'd2033, 32'd1060},
{-32'd408, -32'd1606, -32'd3614, -32'd551},
{-32'd2754, -32'd5554, -32'd2589, -32'd1165},
{-32'd1688, 32'd2652, 32'd6481, 32'd3827},
{32'd8990, -32'd7435, 32'd7993, -32'd51},
{-32'd7988, 32'd3471, -32'd1601, 32'd8233},
{-32'd6434, -32'd2921, -32'd235, -32'd7346},
{32'd1959, -32'd1356, 32'd7947, 32'd3906},
{-32'd1483, 32'd7203, 32'd7890, 32'd797},
{32'd10706, -32'd6668, -32'd5744, 32'd11062},
{32'd2958, -32'd499, -32'd8487, -32'd4999},
{-32'd9072, 32'd5287, -32'd6486, 32'd11235},
{-32'd2950, -32'd3100, -32'd4186, 32'd2610},
{32'd3913, 32'd2741, 32'd3878, 32'd9389},
{32'd5556, -32'd7732, -32'd4817, 32'd1393},
{32'd4640, 32'd1629, -32'd666, 32'd6839},
{-32'd15852, -32'd5783, 32'd916, 32'd609},
{32'd3549, 32'd1453, -32'd1265, 32'd2576},
{-32'd1429, -32'd369, 32'd2875, -32'd5345},
{32'd647, 32'd1955, 32'd5744, 32'd5127},
{-32'd2212, 32'd7069, -32'd5417, -32'd3270},
{-32'd6784, 32'd131, -32'd11863, -32'd3281},
{32'd10360, 32'd4921, -32'd859, -32'd191},
{32'd7084, -32'd2313, 32'd1927, -32'd934},
{-32'd2032, -32'd8301, -32'd9240, -32'd5304},
{32'd2244, 32'd1561, -32'd5612, 32'd6769},
{32'd4565, 32'd5012, 32'd8558, 32'd4621},
{32'd799, -32'd6780, -32'd5358, -32'd1018},
{-32'd1907, 32'd1208, 32'd368, 32'd5779},
{32'd6304, 32'd9470, -32'd5429, -32'd5066},
{-32'd4843, 32'd656, -32'd2807, -32'd6813},
{-32'd4160, -32'd1836, 32'd1083, 32'd8634},
{-32'd6113, -32'd5667, 32'd2249, 32'd5525},
{-32'd5533, 32'd1530, -32'd2876, 32'd3051},
{-32'd1891, 32'd2332, 32'd3826, 32'd3810},
{-32'd7211, -32'd18445, 32'd907, 32'd7843},
{-32'd6918, -32'd2800, 32'd2675, 32'd1427},
{32'd12729, 32'd6654, -32'd3077, -32'd1550},
{-32'd13642, -32'd2776, -32'd2978, 32'd988},
{32'd897, 32'd7443, 32'd490, -32'd2005},
{-32'd8792, 32'd786, -32'd10863, -32'd7510},
{32'd454, 32'd5362, -32'd2498, 32'd3226},
{32'd4354, 32'd6181, 32'd2542, 32'd3926},
{32'd688, -32'd5411, 32'd605, -32'd4975},
{32'd3733, -32'd8494, -32'd4308, -32'd130},
{-32'd788, 32'd5808, 32'd858, 32'd1567},
{-32'd4727, 32'd1227, 32'd5822, -32'd6421},
{-32'd10936, 32'd1365, 32'd5917, -32'd130},
{32'd4354, 32'd1346, -32'd3726, -32'd644},
{-32'd3404, -32'd279, -32'd3259, 32'd599},
{-32'd4913, -32'd7721, -32'd2277, -32'd3031},
{32'd4450, -32'd2920, -32'd3613, -32'd5850},
{-32'd181, -32'd1839, 32'd863, -32'd552},
{32'd12556, -32'd8405, 32'd3194, 32'd5055},
{-32'd13446, -32'd1854, 32'd2988, -32'd8135},
{-32'd824, 32'd2775, -32'd2138, -32'd697},
{-32'd1562, -32'd5599, -32'd5621, -32'd11532},
{-32'd5226, -32'd8313, -32'd3271, 32'd213},
{32'd9103, 32'd9451, 32'd7271, 32'd4403},
{32'd1536, -32'd180, -32'd3934, 32'd5841},
{-32'd5465, -32'd4078, -32'd6816, -32'd4591},
{-32'd4103, 32'd5455, 32'd2561, -32'd6342},
{32'd11822, 32'd1792, -32'd641, -32'd861},
{32'd6656, 32'd15558, 32'd8683, 32'd2667},
{32'd503, 32'd444, 32'd4644, 32'd2108},
{-32'd395, -32'd7859, -32'd4193, 32'd6645},
{-32'd5176, 32'd3434, 32'd7889, 32'd3492},
{-32'd2499, 32'd549, -32'd1843, -32'd6081},
{32'd12107, -32'd1821, 32'd1525, -32'd1168},
{-32'd6920, 32'd3395, -32'd5963, 32'd2485},
{32'd15509, 32'd1312, 32'd11416, -32'd8368},
{32'd4798, 32'd2523, -32'd3459, -32'd8876},
{-32'd2688, 32'd2600, -32'd773, 32'd943},
{32'd8186, 32'd8376, 32'd4097, -32'd3938},
{32'd1976, 32'd4746, 32'd6689, -32'd6202},
{-32'd6600, 32'd2518, -32'd1050, -32'd3415},
{-32'd5284, 32'd6060, -32'd7937, -32'd4290},
{-32'd881, -32'd2473, -32'd6678, 32'd5559},
{-32'd1799, 32'd320, 32'd4918, -32'd230},
{-32'd3209, 32'd5133, 32'd4899, -32'd738},
{32'd7181, 32'd1891, 32'd2568, 32'd873},
{-32'd2889, -32'd5925, -32'd2381, -32'd6874}
},
{{32'd4470, -32'd12178, -32'd1120, 32'd802},
{-32'd7794, -32'd2250, -32'd1883, -32'd1174},
{32'd13608, 32'd237, 32'd8969, -32'd14323},
{32'd8722, 32'd13339, 32'd10474, 32'd4270},
{32'd7622, -32'd509, -32'd821, 32'd7260},
{-32'd3452, 32'd1119, -32'd4661, -32'd6903},
{32'd1081, 32'd6770, 32'd4537, 32'd6142},
{-32'd5245, 32'd1278, 32'd3642, 32'd1278},
{-32'd1701, -32'd3147, 32'd9623, -32'd3532},
{32'd4601, 32'd8780, -32'd1952, 32'd6070},
{-32'd876, -32'd12295, 32'd9877, 32'd7670},
{-32'd7375, 32'd6668, -32'd5029, 32'd8034},
{32'd468, -32'd762, 32'd1881, 32'd4453},
{-32'd99, 32'd1340, -32'd6606, 32'd2843},
{-32'd4165, -32'd5792, 32'd1788, -32'd2443},
{32'd1637, -32'd892, 32'd3223, -32'd634},
{32'd1317, -32'd3047, 32'd10158, 32'd6655},
{-32'd6112, 32'd5433, -32'd9971, -32'd3413},
{32'd5660, 32'd6491, -32'd8353, -32'd3645},
{-32'd4777, 32'd5618, -32'd73, -32'd66},
{32'd3798, -32'd9553, 32'd5127, 32'd7741},
{-32'd675, -32'd2711, 32'd2399, -32'd46},
{32'd3474, -32'd580, 32'd2683, -32'd7986},
{-32'd8528, -32'd2395, -32'd6713, -32'd6230},
{-32'd1869, 32'd4759, 32'd8760, 32'd7936},
{32'd5916, -32'd9406, -32'd2779, 32'd1486},
{-32'd5978, -32'd10711, 32'd3122, 32'd4695},
{-32'd5089, 32'd6703, -32'd5892, -32'd768},
{-32'd6738, 32'd10565, 32'd15868, -32'd7007},
{-32'd5434, -32'd9328, 32'd2544, 32'd3967},
{32'd1139, 32'd3255, 32'd7329, 32'd1210},
{-32'd5088, 32'd835, -32'd5667, -32'd6845},
{32'd11015, 32'd2931, -32'd12191, 32'd2241},
{-32'd3982, -32'd1571, -32'd4616, 32'd4795},
{32'd1925, 32'd8233, 32'd1033, 32'd3956},
{-32'd4098, -32'd2010, 32'd10276, 32'd2842},
{32'd1477, -32'd5051, -32'd9092, -32'd276},
{-32'd4639, -32'd15391, -32'd11274, -32'd5811},
{32'd2004, -32'd7911, -32'd10224, -32'd5198},
{-32'd2663, 32'd5367, 32'd16425, 32'd5873},
{-32'd781, -32'd7429, -32'd4116, -32'd2485},
{-32'd2993, 32'd9362, 32'd14202, 32'd4841},
{-32'd5367, -32'd9990, 32'd9805, 32'd2441},
{-32'd8956, -32'd1524, -32'd2365, -32'd1085},
{32'd2240, -32'd7117, -32'd16830, -32'd2290},
{-32'd3360, -32'd8056, 32'd4488, -32'd1039},
{-32'd6632, 32'd3861, -32'd255, -32'd9481},
{-32'd8770, 32'd5577, -32'd11110, -32'd3872},
{-32'd1769, 32'd1972, 32'd579, 32'd8290},
{-32'd3550, -32'd1834, -32'd5917, -32'd1198},
{32'd2284, -32'd5595, -32'd3866, -32'd345},
{-32'd5552, 32'd4686, -32'd10464, 32'd6573},
{32'd2084, 32'd5996, -32'd2766, -32'd13483},
{-32'd2354, -32'd11797, -32'd1974, 32'd2283},
{32'd6713, -32'd6600, 32'd2501, -32'd4749},
{-32'd1350, -32'd2610, -32'd6922, -32'd34},
{32'd14688, 32'd9655, -32'd10017, -32'd652},
{-32'd541, -32'd5848, -32'd10294, 32'd224},
{-32'd3894, -32'd11960, -32'd261, -32'd473},
{-32'd8080, -32'd775, 32'd10154, 32'd1932},
{32'd3110, -32'd2824, -32'd3237, 32'd7890},
{32'd1171, 32'd410, 32'd7976, -32'd1747},
{-32'd5176, 32'd3923, 32'd4496, -32'd317},
{-32'd540, -32'd3382, 32'd5782, 32'd8192},
{-32'd2431, -32'd12739, -32'd4587, -32'd5903},
{32'd1375, 32'd9158, 32'd8069, 32'd8264},
{-32'd12321, -32'd408, 32'd8084, 32'd4243},
{-32'd3120, 32'd4569, -32'd3402, -32'd1020},
{-32'd3096, -32'd10167, -32'd2904, -32'd3399},
{32'd1689, 32'd9191, 32'd13853, 32'd644},
{32'd2202, -32'd4688, 32'd126, -32'd8578},
{-32'd2599, -32'd2754, 32'd14282, -32'd5527},
{32'd2928, -32'd13941, 32'd2243, -32'd16693},
{32'd3022, -32'd9797, 32'd4657, 32'd10473},
{32'd11800, -32'd8504, -32'd4306, -32'd3273},
{32'd2375, -32'd480, 32'd7166, -32'd3736},
{32'd3073, 32'd1242, -32'd6422, -32'd2598},
{-32'd1429, -32'd4286, -32'd2854, 32'd8003},
{32'd6147, 32'd4050, 32'd12167, 32'd5892},
{32'd7006, 32'd1830, -32'd2551, -32'd3354},
{32'd9214, -32'd5193, -32'd7531, 32'd2251},
{32'd2362, -32'd3679, 32'd137, 32'd7391},
{32'd3309, -32'd12056, -32'd2206, 32'd2745},
{32'd7471, -32'd7840, 32'd3178, -32'd5656},
{-32'd731, -32'd7587, -32'd6593, 32'd11262},
{32'd4191, -32'd5994, 32'd4135, -32'd6820},
{32'd10484, -32'd925, 32'd4061, -32'd8537},
{-32'd3162, 32'd1453, -32'd3046, -32'd1938},
{32'd1746, -32'd677, -32'd8147, -32'd4665},
{32'd2144, 32'd2548, -32'd5102, -32'd18213},
{-32'd6, -32'd2992, 32'd4823, 32'd6398},
{-32'd6512, -32'd9763, 32'd4557, 32'd3888},
{-32'd6716, 32'd9866, -32'd1693, 32'd3997},
{32'd3749, 32'd6475, 32'd621, 32'd6157},
{32'd584, 32'd1309, 32'd2459, -32'd1951},
{32'd2625, -32'd6255, 32'd957, -32'd4812},
{-32'd628, -32'd2449, -32'd1424, 32'd5697},
{32'd3796, 32'd2443, 32'd3938, -32'd8756},
{-32'd6213, 32'd7051, 32'd747, -32'd386},
{32'd3029, 32'd4265, 32'd6205, -32'd2052},
{-32'd6892, 32'd7843, 32'd1373, -32'd6268},
{32'd2030, 32'd5618, 32'd11073, 32'd3437},
{32'd8145, 32'd2535, -32'd8569, 32'd5402},
{-32'd3407, 32'd1055, 32'd8012, -32'd3980},
{32'd4430, -32'd6685, 32'd2617, -32'd694},
{32'd192, 32'd11518, 32'd7848, 32'd14121},
{-32'd7730, -32'd3458, -32'd1392, -32'd5774},
{32'd5167, 32'd865, 32'd14155, -32'd1132},
{32'd114, 32'd8909, -32'd165, -32'd1390},
{32'd3375, -32'd676, 32'd3381, -32'd3308},
{32'd3972, -32'd3380, -32'd1024, 32'd4145},
{32'd1129, -32'd4381, -32'd2943, -32'd4624},
{-32'd814, 32'd2565, 32'd3957, 32'd8378},
{-32'd7562, 32'd11558, -32'd4083, 32'd15176},
{-32'd3287, -32'd3315, 32'd3680, -32'd8238},
{32'd2171, -32'd3186, 32'd2794, -32'd2017},
{-32'd6825, 32'd9489, 32'd13276, 32'd10293},
{-32'd2375, -32'd1031, 32'd4711, -32'd3142},
{-32'd7361, 32'd4496, -32'd3131, 32'd13208},
{32'd1235, 32'd11741, 32'd8511, 32'd6844},
{-32'd191, -32'd1779, 32'd6413, -32'd2146},
{32'd6965, -32'd1821, -32'd1791, -32'd5319},
{-32'd3676, 32'd4581, -32'd136, 32'd1058},
{32'd1532, 32'd4694, 32'd6133, -32'd5420},
{-32'd3141, 32'd5269, -32'd3763, 32'd2928},
{-32'd917, 32'd8747, 32'd8072, -32'd5722},
{32'd6411, -32'd6636, -32'd4933, 32'd8904},
{-32'd3972, -32'd3680, 32'd7355, -32'd6227},
{32'd730, -32'd2048, 32'd6170, -32'd13161},
{32'd4006, -32'd17279, 32'd4134, 32'd7182},
{32'd5607, -32'd1598, -32'd11013, 32'd1030},
{-32'd4393, -32'd3779, -32'd9255, -32'd5700},
{-32'd2805, -32'd8009, 32'd7150, 32'd1443},
{-32'd1389, -32'd4367, -32'd2426, -32'd5099},
{32'd2553, 32'd23122, 32'd6746, -32'd3879},
{32'd8973, 32'd2580, 32'd5664, 32'd10457},
{-32'd4276, 32'd6916, -32'd2153, 32'd12998},
{-32'd2398, 32'd121, -32'd5760, 32'd172},
{-32'd1935, 32'd13387, -32'd4013, 32'd4976},
{32'd6179, -32'd15579, -32'd4442, 32'd5416},
{32'd5672, -32'd10053, -32'd9011, 32'd2346},
{-32'd1105, -32'd3023, -32'd1327, -32'd1951},
{-32'd6360, 32'd5722, 32'd4077, 32'd7998},
{32'd9713, 32'd626, -32'd1121, -32'd3655},
{-32'd152, 32'd2161, 32'd4863, 32'd1531},
{32'd6436, 32'd588, -32'd5728, 32'd11881},
{-32'd6851, -32'd11253, -32'd4980, 32'd7479},
{-32'd2269, -32'd3131, -32'd2127, 32'd1193},
{32'd3632, 32'd18736, -32'd5027, 32'd1465},
{32'd158, 32'd1611, -32'd14858, 32'd4287},
{-32'd4333, -32'd11084, -32'd2630, -32'd136},
{32'd359, 32'd7679, -32'd1598, 32'd856},
{-32'd10414, 32'd12971, 32'd2377, 32'd6722},
{32'd4769, -32'd10801, 32'd4940, 32'd5013},
{-32'd9961, -32'd6981, 32'd3774, -32'd2494},
{32'd9050, 32'd683, -32'd3820, 32'd900},
{32'd3323, 32'd3058, -32'd5026, -32'd1402},
{-32'd4639, -32'd1937, 32'd14462, -32'd8650},
{-32'd5128, -32'd9229, -32'd4501, -32'd2825},
{32'd397, -32'd12898, -32'd3887, 32'd1191},
{-32'd3406, -32'd4677, 32'd5056, -32'd12720},
{-32'd4032, 32'd3561, -32'd5954, -32'd5320},
{-32'd14494, 32'd0, 32'd1163, 32'd107},
{32'd6129, 32'd12772, 32'd8351, 32'd3706},
{32'd4928, 32'd1889, 32'd9725, -32'd616},
{-32'd3132, -32'd7415, -32'd4925, -32'd9013},
{-32'd2106, 32'd8176, 32'd8750, -32'd9159},
{32'd5342, -32'd7549, -32'd3823, -32'd10128},
{32'd3021, -32'd12303, 32'd1141, -32'd5885},
{32'd1741, -32'd2802, 32'd10463, -32'd1023},
{-32'd8148, -32'd11426, -32'd1175, 32'd6424},
{-32'd9697, -32'd64, -32'd2915, 32'd7980},
{32'd4940, 32'd9044, 32'd7286, 32'd3037},
{-32'd4206, -32'd3023, 32'd9202, 32'd2622},
{32'd3113, 32'd11344, -32'd5530, 32'd10310},
{32'd4204, -32'd4168, 32'd679, -32'd6926},
{32'd10747, 32'd5976, 32'd203, -32'd1767},
{-32'd4525, 32'd8208, 32'd1414, 32'd1617},
{-32'd8255, 32'd13175, 32'd3371, 32'd11944},
{-32'd1711, -32'd3924, -32'd11809, -32'd6542},
{-32'd8686, -32'd6432, 32'd7656, 32'd2953},
{32'd1885, -32'd8599, -32'd2805, -32'd3571},
{-32'd4396, 32'd2175, -32'd228, -32'd6157},
{-32'd11036, -32'd7774, -32'd31, 32'd7711},
{-32'd3389, 32'd4548, 32'd4282, -32'd1289},
{32'd6407, -32'd287, -32'd1530, 32'd3364},
{32'd4023, 32'd12055, 32'd17776, 32'd2279},
{-32'd10269, 32'd7118, 32'd6894, -32'd2218},
{32'd3112, 32'd5801, -32'd2965, -32'd6654},
{32'd7708, -32'd9208, -32'd914, -32'd447},
{-32'd3993, 32'd65, 32'd397, -32'd1834},
{32'd1959, 32'd240, 32'd1749, -32'd10003},
{-32'd11962, 32'd3463, 32'd10411, -32'd4835},
{32'd4786, 32'd9852, -32'd16473, -32'd4784},
{-32'd2435, 32'd5749, -32'd7114, -32'd6949},
{-32'd5009, 32'd979, 32'd2419, 32'd4995},
{-32'd10668, 32'd8809, -32'd4544, -32'd761},
{32'd9699, -32'd5693, -32'd1043, 32'd7460},
{32'd5713, -32'd5297, -32'd10140, 32'd8625},
{-32'd3221, -32'd8428, 32'd7237, 32'd3165},
{-32'd6048, -32'd8256, -32'd4134, -32'd2620},
{-32'd7109, -32'd6655, 32'd10830, 32'd13967},
{-32'd2233, 32'd1446, -32'd8152, 32'd16566},
{32'd1419, 32'd8980, 32'd3765, 32'd2547},
{-32'd4403, 32'd2180, -32'd3051, -32'd7543},
{-32'd2013, 32'd3742, 32'd4688, -32'd3804},
{-32'd2472, 32'd8376, 32'd3130, 32'd3517},
{-32'd3202, -32'd11807, -32'd10328, -32'd838},
{32'd6615, 32'd21158, 32'd4034, -32'd1909},
{32'd4198, 32'd426, 32'd5050, 32'd2044},
{32'd5007, -32'd4801, -32'd5890, -32'd3741},
{32'd206, -32'd12768, -32'd5800, 32'd1825},
{32'd6361, 32'd1780, -32'd3632, -32'd6788},
{-32'd7206, -32'd7766, -32'd6222, 32'd371},
{32'd4359, -32'd15977, -32'd3822, 32'd9044},
{-32'd4892, 32'd11220, -32'd2225, -32'd4},
{-32'd9977, -32'd124, -32'd2365, 32'd5469},
{32'd6553, -32'd6184, -32'd3383, -32'd8858},
{32'd2250, -32'd2021, -32'd158, 32'd10113},
{-32'd6622, 32'd6778, -32'd6450, 32'd1519},
{-32'd8517, -32'd641, -32'd4721, -32'd1630},
{-32'd8293, 32'd4789, 32'd5442, 32'd5905},
{32'd1542, 32'd5240, 32'd6948, -32'd4210},
{-32'd4047, -32'd3656, -32'd1854, 32'd4605},
{32'd7392, -32'd1535, -32'd1772, -32'd3510},
{32'd3816, 32'd4867, -32'd5034, 32'd3186},
{-32'd5480, 32'd2178, -32'd9081, 32'd1543},
{-32'd2025, -32'd3920, 32'd11713, -32'd11081},
{-32'd4714, 32'd12115, -32'd2394, 32'd5254},
{32'd5218, 32'd98, 32'd6702, -32'd4197},
{-32'd3727, -32'd2256, 32'd3903, 32'd3630},
{-32'd8343, 32'd6116, 32'd14212, 32'd9877},
{32'd10686, -32'd89, 32'd3117, -32'd6213},
{32'd7668, 32'd8307, 32'd4779, -32'd2904},
{32'd286, -32'd4197, -32'd12615, -32'd13935},
{-32'd7682, 32'd370, -32'd8915, -32'd4608},
{32'd218, 32'd330, -32'd14968, 32'd178},
{32'd7678, -32'd10642, -32'd6038, -32'd5087},
{32'd3715, -32'd4205, 32'd8818, -32'd2715},
{-32'd445, -32'd713, 32'd7942, -32'd1853},
{32'd1104, 32'd2315, 32'd8588, 32'd9874},
{-32'd3303, -32'd10, -32'd2430, 32'd8648},
{32'd73, -32'd8360, 32'd6498, -32'd5390},
{32'd9694, -32'd7513, -32'd2616, -32'd6773},
{32'd7119, 32'd5867, -32'd2279, 32'd11560},
{32'd3082, -32'd3451, -32'd7197, -32'd34},
{-32'd2704, -32'd8258, -32'd11725, -32'd6771},
{-32'd1121, 32'd5392, 32'd3293, -32'd11685},
{32'd5811, 32'd6188, -32'd210, -32'd5390},
{32'd3587, -32'd6932, -32'd2117, 32'd495},
{-32'd4110, 32'd1117, -32'd1012, -32'd3236},
{32'd2982, 32'd11358, -32'd3366, 32'd293},
{-32'd2355, -32'd4509, -32'd2995, -32'd3818},
{-32'd1376, 32'd4519, -32'd11417, 32'd3852},
{-32'd143, -32'd5591, -32'd6228, 32'd435},
{32'd2980, 32'd3002, 32'd1473, -32'd500},
{-32'd8930, 32'd4794, -32'd8784, 32'd6663},
{32'd6671, 32'd4090, -32'd3614, 32'd2679},
{-32'd9902, -32'd4749, 32'd411, 32'd3605},
{-32'd3961, 32'd176, -32'd11096, -32'd518},
{-32'd4432, 32'd20494, 32'd7006, 32'd5450},
{32'd5608, 32'd6963, -32'd7698, -32'd986},
{32'd348, -32'd8029, -32'd4339, -32'd2779},
{-32'd36, -32'd1967, 32'd953, 32'd712},
{-32'd386, 32'd1198, 32'd10165, -32'd4645},
{32'd6003, -32'd2779, -32'd9482, 32'd3952},
{32'd11861, 32'd8978, -32'd1741, 32'd77},
{-32'd1723, -32'd2232, 32'd9001, -32'd4453},
{-32'd4931, 32'd2495, 32'd8772, 32'd6759},
{-32'd8330, 32'd908, -32'd2401, -32'd1136},
{32'd3888, -32'd2376, -32'd5627, -32'd8981},
{32'd2256, -32'd3509, 32'd6852, -32'd12291},
{-32'd2408, 32'd828, -32'd5124, -32'd8642},
{-32'd11351, 32'd1326, 32'd11217, -32'd8350},
{32'd2777, -32'd7791, -32'd141, -32'd2415},
{-32'd3248, -32'd9767, -32'd2255, -32'd1736},
{32'd6794, 32'd11393, 32'd1690, 32'd6855},
{-32'd10073, -32'd4468, 32'd10143, 32'd2841},
{32'd863, -32'd1629, -32'd4699, -32'd4728},
{32'd6443, 32'd7463, 32'd1008, -32'd6330},
{32'd4857, 32'd1590, -32'd982, -32'd2565},
{-32'd2774, -32'd898, 32'd9563, 32'd6305},
{32'd8529, -32'd6761, 32'd11692, -32'd741},
{32'd7086, 32'd3793, -32'd136, 32'd3543},
{32'd8648, 32'd1039, 32'd5124, 32'd5498},
{-32'd5199, -32'd16100, -32'd9700, -32'd13070},
{-32'd4768, 32'd9110, -32'd2731, -32'd1590},
{-32'd2049, -32'd15581, -32'd3037, -32'd5125},
{-32'd5159, 32'd1061, 32'd9684, 32'd1027},
{32'd4468, -32'd1327, -32'd13516, -32'd7950},
{32'd4979, 32'd13923, 32'd3381, 32'd5222},
{32'd11981, 32'd10189, 32'd8934, -32'd2680},
{32'd2355, -32'd6236, -32'd5946, -32'd6733},
{32'd12457, 32'd15, -32'd5184, -32'd753},
{-32'd675, -32'd1459, -32'd5577, -32'd8059},
{-32'd8159, -32'd9871, -32'd8561, 32'd634},
{32'd1045, -32'd4369, 32'd2768, 32'd1382},
{32'd2741, 32'd12464, 32'd7934, -32'd644},
{32'd10921, 32'd16179, 32'd797, -32'd3181},
{32'd1762, -32'd20244, -32'd10122, 32'd5153}
},
{{-32'd3966, -32'd4336, 32'd5236, 32'd2580},
{-32'd12996, -32'd5454, -32'd4062, 32'd4605},
{-32'd5340, 32'd9337, 32'd127, -32'd9244},
{32'd12410, -32'd4318, 32'd1149, 32'd11881},
{-32'd3426, 32'd6899, 32'd8585, -32'd3666},
{32'd2694, 32'd1116, -32'd8820, 32'd2716},
{32'd1024, -32'd2259, 32'd10053, -32'd1388},
{32'd6397, -32'd13835, -32'd5932, -32'd11646},
{32'd369, 32'd10565, -32'd273, 32'd1227},
{32'd6950, 32'd4705, 32'd2772, 32'd12644},
{-32'd3049, -32'd4308, -32'd7438, -32'd3478},
{32'd3604, 32'd5116, -32'd9809, -32'd3773},
{32'd7852, -32'd5659, 32'd5099, 32'd11342},
{32'd2087, -32'd15580, -32'd1637, 32'd122},
{-32'd4618, -32'd12448, -32'd7779, -32'd2089},
{32'd1903, -32'd50, -32'd1690, -32'd2879},
{32'd8913, -32'd3166, -32'd768, -32'd360},
{-32'd6541, -32'd1265, 32'd578, -32'd1464},
{-32'd2598, -32'd10420, 32'd3763, -32'd3561},
{-32'd3539, 32'd2218, -32'd9870, -32'd382},
{32'd4448, 32'd9656, -32'd315, 32'd6049},
{-32'd220, 32'd929, -32'd5635, 32'd1887},
{-32'd3941, -32'd4603, -32'd1512, 32'd6563},
{-32'd1972, -32'd1103, -32'd3067, -32'd3521},
{32'd2072, 32'd3133, 32'd703, 32'd2649},
{32'd3143, -32'd6417, -32'd3092, -32'd8667},
{-32'd1310, 32'd1875, 32'd9434, 32'd8497},
{32'd9607, 32'd4617, -32'd148, -32'd6545},
{32'd4368, -32'd2918, 32'd5741, -32'd4687},
{-32'd1249, -32'd6300, 32'd6026, 32'd858},
{-32'd1601, -32'd2826, -32'd12518, -32'd1469},
{-32'd8900, -32'd10516, 32'd1135, -32'd8828},
{32'd4920, 32'd3555, 32'd12472, 32'd4640},
{32'd1421, -32'd2797, -32'd2632, -32'd5289},
{32'd9458, 32'd14816, 32'd4611, 32'd6935},
{-32'd7107, 32'd4069, 32'd10435, -32'd3437},
{32'd4207, -32'd7943, 32'd3603, -32'd10271},
{32'd4585, -32'd11715, 32'd568, -32'd4297},
{32'd969, -32'd12796, -32'd1825, 32'd5991},
{32'd2126, 32'd4338, 32'd3102, -32'd3038},
{32'd8218, -32'd509, -32'd10218, -32'd2710},
{32'd722, 32'd9499, 32'd8264, 32'd164},
{-32'd5252, -32'd4293, -32'd7140, -32'd5601},
{-32'd765, -32'd17576, -32'd3826, 32'd1232},
{-32'd4621, -32'd7673, 32'd2151, -32'd6739},
{-32'd3315, 32'd52, -32'd7381, 32'd7491},
{-32'd11958, -32'd1220, 32'd1939, -32'd5107},
{-32'd907, -32'd6592, -32'd4813, -32'd8976},
{32'd1913, 32'd5819, 32'd6586, 32'd1484},
{-32'd3997, -32'd4437, 32'd4885, -32'd3853},
{-32'd6155, 32'd1673, 32'd7206, -32'd5345},
{32'd2926, 32'd4894, -32'd728, -32'd2489},
{-32'd5073, 32'd6112, -32'd1480, -32'd1311},
{-32'd8901, -32'd1622, -32'd5405, 32'd2797},
{32'd1271, 32'd4252, 32'd124, 32'd7994},
{-32'd577, -32'd10346, -32'd2082, 32'd6032},
{-32'd191, -32'd2870, -32'd371, -32'd1306},
{-32'd14035, -32'd5258, -32'd6498, -32'd12420},
{-32'd1707, -32'd2190, -32'd7196, -32'd9572},
{-32'd3986, 32'd9880, -32'd1770, -32'd3108},
{-32'd5726, 32'd4924, 32'd7500, 32'd9560},
{32'd5852, -32'd4828, 32'd15347, -32'd5299},
{-32'd14606, -32'd9670, -32'd1304, -32'd13936},
{-32'd8713, 32'd8371, 32'd7883, 32'd2950},
{-32'd491, 32'd3231, 32'd1128, 32'd6999},
{32'd1690, 32'd3875, 32'd9747, 32'd6637},
{32'd2863, -32'd10202, -32'd11834, 32'd8089},
{-32'd12697, -32'd386, -32'd6581, 32'd2385},
{-32'd7067, -32'd4997, -32'd3757, -32'd1086},
{32'd3127, 32'd1530, 32'd294, 32'd2995},
{-32'd5570, 32'd5304, -32'd1286, -32'd6770},
{-32'd3772, 32'd6474, 32'd12198, -32'd964},
{-32'd7129, 32'd4238, 32'd2810, -32'd10883},
{32'd7491, 32'd2865, -32'd2153, 32'd5804},
{32'd10691, 32'd368, 32'd3509, 32'd6485},
{-32'd2264, -32'd3565, 32'd10632, 32'd5289},
{-32'd8262, -32'd5820, -32'd9128, -32'd321},
{32'd9554, 32'd373, -32'd3210, -32'd8765},
{32'd1642, 32'd204, 32'd12659, 32'd1354},
{-32'd3284, 32'd1501, -32'd2584, -32'd1123},
{32'd3369, 32'd950, 32'd11054, -32'd13301},
{-32'd3047, -32'd6575, 32'd14343, 32'd11675},
{32'd327, 32'd16, 32'd7184, 32'd1329},
{-32'd243, 32'd1208, -32'd1154, -32'd478},
{-32'd9138, -32'd4816, -32'd2666, -32'd5500},
{-32'd5606, 32'd3468, 32'd2619, -32'd3791},
{32'd1823, 32'd4219, -32'd3203, -32'd9052},
{-32'd1860, 32'd3936, 32'd5436, -32'd17214},
{-32'd10294, 32'd1590, 32'd2305, 32'd777},
{-32'd4343, 32'd2345, 32'd1274, -32'd2180},
{-32'd5759, -32'd8162, -32'd3184, 32'd1510},
{-32'd629, -32'd3837, 32'd1569, -32'd4718},
{32'd2148, -32'd2033, -32'd588, -32'd1234},
{32'd8139, 32'd2219, 32'd3008, 32'd5815},
{-32'd5570, -32'd3781, 32'd6387, -32'd7870},
{-32'd3483, -32'd11834, -32'd5029, -32'd6641},
{32'd5851, 32'd3804, 32'd1470, -32'd979},
{32'd5917, 32'd5958, 32'd1868, 32'd1737},
{32'd6705, 32'd520, 32'd10340, -32'd4285},
{32'd6539, 32'd1667, -32'd7086, 32'd469},
{-32'd7542, -32'd2195, -32'd8776, 32'd3442},
{32'd1839, -32'd8315, 32'd7805, -32'd3139},
{-32'd6726, -32'd2726, 32'd859, 32'd8724},
{32'd7474, 32'd9594, -32'd4517, 32'd3233},
{32'd9435, 32'd11204, 32'd10839, 32'd2412},
{-32'd8036, -32'd577, -32'd6089, 32'd5141},
{-32'd2380, 32'd3491, -32'd337, 32'd2653},
{-32'd2784, 32'd2625, 32'd3213, 32'd548},
{32'd4247, -32'd1913, 32'd1851, 32'd18011},
{-32'd9327, 32'd3166, -32'd2461, -32'd2315},
{32'd2787, -32'd4122, 32'd7553, -32'd6978},
{-32'd2478, 32'd6831, 32'd2468, -32'd3232},
{-32'd592, 32'd5900, 32'd4998, 32'd5802},
{-32'd1293, 32'd6747, -32'd2954, 32'd1350},
{-32'd7783, -32'd6256, -32'd3934, 32'd5063},
{-32'd474, 32'd5382, 32'd5736, 32'd5687},
{32'd7591, 32'd4954, 32'd1586, -32'd4836},
{-32'd1903, -32'd4485, 32'd1664, 32'd2886},
{32'd8871, -32'd8341, 32'd12186, -32'd969},
{32'd9789, 32'd11675, 32'd7762, 32'd10058},
{-32'd4264, -32'd7434, -32'd2873, 32'd2138},
{32'd8330, 32'd2010, -32'd3255, 32'd8601},
{-32'd1738, 32'd12631, -32'd5178, 32'd7259},
{32'd6009, -32'd8488, -32'd11700, -32'd5250},
{-32'd6829, 32'd5253, 32'd10362, -32'd527},
{32'd3258, -32'd9375, -32'd1799, 32'd11134},
{-32'd2370, 32'd153, -32'd1847, -32'd3405},
{32'd150, -32'd5279, -32'd2038, -32'd10687},
{-32'd1473, -32'd2581, -32'd15323, 32'd1641},
{32'd1958, 32'd3431, 32'd2081, -32'd1984},
{32'd4030, 32'd15964, 32'd9779, 32'd3665},
{-32'd14750, -32'd12059, 32'd3932, -32'd5648},
{32'd1114, -32'd10919, -32'd8798, -32'd12808},
{32'd1559, 32'd2014, 32'd4749, -32'd4523},
{-32'd4780, 32'd7565, -32'd1613, -32'd1654},
{32'd8082, -32'd5274, 32'd7320, -32'd5622},
{-32'd13791, 32'd4075, 32'd8527, 32'd439},
{32'd3484, -32'd9022, -32'd13708, 32'd10285},
{-32'd5529, 32'd1565, -32'd685, -32'd207},
{32'd158, -32'd5874, -32'd9501, -32'd9741},
{32'd3438, -32'd3335, -32'd2319, 32'd1118},
{32'd92, 32'd196, -32'd5609, -32'd21631},
{-32'd3260, -32'd8506, 32'd2349, -32'd885},
{32'd3963, 32'd5250, 32'd2284, -32'd3986},
{-32'd246, 32'd6977, -32'd3236, 32'd1941},
{32'd6033, -32'd984, 32'd6310, 32'd4777},
{32'd6198, -32'd1225, -32'd4485, -32'd8565},
{32'd4178, -32'd4863, -32'd3283, 32'd1034},
{32'd7336, 32'd1383, 32'd5731, 32'd381},
{-32'd542, -32'd4241, -32'd7479, -32'd818},
{-32'd4205, -32'd12446, -32'd4426, -32'd12154},
{32'd3472, -32'd6942, -32'd2133, 32'd7547},
{32'd2600, -32'd4522, 32'd8082, 32'd3156},
{-32'd4919, -32'd2278, -32'd3462, 32'd4462},
{-32'd20087, 32'd767, -32'd6921, -32'd12746},
{32'd1509, -32'd12141, -32'd2366, 32'd1839},
{-32'd3913, 32'd14817, 32'd8760, -32'd800},
{-32'd549, 32'd3119, -32'd1320, 32'd4229},
{32'd3210, 32'd3669, 32'd2210, 32'd2593},
{-32'd6747, -32'd354, 32'd4957, -32'd12668},
{32'd5664, 32'd1913, -32'd3824, -32'd427},
{32'd3058, -32'd9554, 32'd992, 32'd4534},
{-32'd1894, 32'd10297, -32'd2660, -32'd12520},
{32'd4342, 32'd2552, -32'd1211, -32'd615},
{32'd1913, 32'd7944, 32'd796, 32'd9864},
{-32'd341, -32'd87, -32'd133, 32'd6090},
{-32'd2231, -32'd6230, -32'd2158, -32'd2686},
{-32'd5786, -32'd6638, -32'd5606, -32'd7433},
{-32'd3948, 32'd2806, 32'd105, -32'd4735},
{-32'd4126, 32'd14, 32'd1171, -32'd6036},
{32'd3924, -32'd2387, -32'd8769, 32'd812},
{-32'd10266, -32'd5806, -32'd8390, 32'd4073},
{32'd8040, 32'd6153, -32'd570, 32'd4886},
{32'd2022, -32'd5721, -32'd1479, -32'd9928},
{32'd9979, -32'd3977, 32'd7392, 32'd9538},
{-32'd1788, -32'd2062, 32'd554, 32'd2472},
{32'd5221, -32'd809, -32'd1150, 32'd3589},
{32'd687, -32'd1504, 32'd9620, 32'd2435},
{32'd8303, -32'd9790, 32'd2105, 32'd1936},
{-32'd1973, -32'd8718, -32'd6339, -32'd2825},
{32'd2037, 32'd1852, 32'd2129, -32'd6052},
{-32'd6147, -32'd9158, -32'd1741, -32'd7148},
{-32'd6209, -32'd9218, -32'd8210, 32'd1332},
{-32'd5378, -32'd677, 32'd1582, 32'd2868},
{-32'd2221, -32'd3739, -32'd2972, 32'd10334},
{32'd7168, 32'd8412, -32'd2637, 32'd4485},
{32'd4606, -32'd1209, -32'd794, 32'd2009},
{32'd4555, -32'd1727, 32'd5298, 32'd10944},
{32'd5889, 32'd1019, 32'd17758, 32'd1104},
{-32'd5279, -32'd1480, -32'd3861, 32'd3613},
{32'd2151, 32'd4899, 32'd7708, -32'd3168},
{-32'd1435, -32'd12131, -32'd2218, -32'd8907},
{-32'd2112, -32'd3892, -32'd594, 32'd6644},
{-32'd3544, -32'd5861, 32'd4672, 32'd2006},
{32'd5930, 32'd1207, 32'd1617, 32'd7664},
{32'd3070, 32'd716, 32'd1989, 32'd3020},
{-32'd9566, -32'd2988, -32'd1112, -32'd4314},
{32'd7701, 32'd10056, 32'd6152, 32'd13108},
{-32'd3089, -32'd4718, 32'd2711, -32'd2811},
{-32'd6542, -32'd2048, -32'd4691, 32'd3707},
{-32'd9261, -32'd11425, -32'd6705, -32'd6310},
{32'd5909, -32'd3359, 32'd2572, -32'd682},
{-32'd1295, 32'd3966, 32'd4821, -32'd3689},
{32'd11460, -32'd5975, -32'd2986, 32'd9693},
{-32'd11097, -32'd4832, -32'd8764, -32'd2031},
{32'd6671, -32'd4803, 32'd5546, 32'd617},
{32'd15131, 32'd6230, -32'd7059, 32'd4565},
{-32'd5706, -32'd12663, -32'd11091, 32'd7602},
{-32'd817, -32'd5680, 32'd2811, -32'd12301},
{-32'd2342, 32'd6405, -32'd5411, -32'd3305},
{-32'd7105, -32'd772, -32'd5087, -32'd277},
{-32'd4307, 32'd7297, 32'd6775, 32'd4965},
{-32'd7621, 32'd1284, 32'd5072, 32'd3511},
{32'd7247, -32'd8275, 32'd9078, 32'd16467},
{-32'd9825, -32'd7896, -32'd9431, -32'd7095},
{-32'd3375, 32'd1513, -32'd6541, -32'd5923},
{-32'd1215, 32'd2713, 32'd1127, 32'd4072},
{32'd7873, -32'd4364, -32'd1797, 32'd3029},
{32'd9145, 32'd4071, 32'd3376, 32'd9878},
{32'd12257, -32'd5031, 32'd7217, 32'd5107},
{-32'd5450, -32'd14287, -32'd1254, 32'd1814},
{32'd7903, 32'd14216, 32'd5587, 32'd1571},
{32'd5422, 32'd664, 32'd19139, -32'd1856},
{-32'd785, 32'd11221, 32'd5310, -32'd1569},
{-32'd4941, 32'd5229, 32'd1421, -32'd696},
{32'd4104, -32'd956, 32'd11197, 32'd2136},
{32'd2111, -32'd1834, -32'd2267, 32'd4674},
{-32'd18923, 32'd174, 32'd3403, -32'd8429},
{32'd8617, -32'd2667, 32'd418, -32'd9952},
{-32'd8180, -32'd2368, -32'd348, 32'd11346},
{-32'd7852, 32'd6729, -32'd1052, -32'd7340},
{32'd4075, -32'd2585, 32'd1953, -32'd3064},
{32'd256, 32'd10810, 32'd7702, 32'd4188},
{-32'd2682, 32'd4613, 32'd1230, -32'd9690},
{-32'd834, -32'd8968, -32'd842, -32'd659},
{-32'd8158, -32'd8107, -32'd8500, -32'd3196},
{32'd4126, 32'd2735, -32'd5081, 32'd2692},
{32'd9575, -32'd20, 32'd12788, 32'd2347},
{32'd4589, 32'd49, 32'd4659, 32'd137},
{-32'd755, 32'd7346, -32'd855, -32'd4666},
{-32'd8639, 32'd6032, 32'd8496, -32'd5083},
{-32'd3477, 32'd3214, -32'd14214, -32'd5709},
{-32'd2265, -32'd8101, -32'd3907, -32'd8283},
{32'd9538, -32'd3503, -32'd1380, 32'd12492},
{32'd9052, 32'd9096, 32'd3339, 32'd13784},
{-32'd696, -32'd3626, -32'd1053, 32'd4578},
{-32'd1967, 32'd1944, 32'd4599, -32'd5671},
{-32'd7345, 32'd7144, -32'd4964, 32'd6429},
{32'd2001, 32'd1332, -32'd5008, 32'd1940},
{32'd6466, -32'd1780, 32'd9273, 32'd10107},
{-32'd4627, -32'd2797, 32'd4840, 32'd11278},
{-32'd3297, 32'd5848, 32'd1155, -32'd7421},
{32'd1243, -32'd3192, -32'd6336, -32'd2538},
{32'd4285, 32'd2309, 32'd7683, 32'd14361},
{32'd15, 32'd899, 32'd3891, -32'd1054},
{32'd755, -32'd3633, -32'd5754, -32'd3233},
{32'd4754, 32'd2988, -32'd6035, 32'd2619},
{32'd14139, -32'd887, 32'd5161, 32'd1210},
{-32'd1832, -32'd2409, -32'd15482, -32'd9011},
{32'd2980, 32'd5676, 32'd6539, 32'd4977},
{32'd1240, 32'd2510, 32'd1471, 32'd2550},
{-32'd3604, -32'd5452, -32'd2894, -32'd1662},
{-32'd3483, -32'd9622, -32'd9803, -32'd4858},
{-32'd2779, -32'd674, 32'd8980, 32'd660},
{32'd1995, 32'd4678, 32'd1803, -32'd1721},
{-32'd5284, -32'd3431, -32'd114, -32'd1715},
{32'd503, 32'd599, 32'd13114, 32'd3023},
{-32'd9539, 32'd3690, -32'd1225, -32'd6230},
{-32'd3345, -32'd5099, -32'd1537, -32'd5075},
{-32'd5771, 32'd5170, -32'd146, -32'd5490},
{32'd1948, 32'd3969, 32'd1428, 32'd9228},
{32'd7749, 32'd7805, -32'd694, 32'd3048},
{-32'd4788, -32'd3890, 32'd1543, -32'd2967},
{-32'd785, 32'd9538, -32'd5345, -32'd2381},
{32'd2083, -32'd3558, -32'd160, 32'd10583},
{-32'd9861, -32'd479, 32'd8109, -32'd5037},
{32'd6260, 32'd9229, 32'd5811, 32'd13200},
{32'd5211, 32'd6951, 32'd2145, 32'd4404},
{-32'd2839, -32'd3632, -32'd6552, -32'd4277},
{-32'd1433, -32'd1537, -32'd6174, 32'd1713},
{32'd4642, 32'd534, 32'd1642, 32'd7246},
{32'd1778, 32'd7715, -32'd4730, 32'd5020},
{32'd7591, 32'd1399, 32'd6102, -32'd8454},
{32'd638, 32'd7947, -32'd2655, 32'd10245},
{-32'd198, -32'd2588, -32'd2160, -32'd7977},
{-32'd2345, -32'd11087, -32'd15888, -32'd12247},
{32'd281, -32'd468, 32'd2118, 32'd5220},
{-32'd3388, 32'd9648, 32'd1319, 32'd5837},
{-32'd6410, 32'd569, -32'd7944, -32'd8825},
{-32'd2888, -32'd3318, -32'd13011, 32'd412},
{32'd8293, -32'd227, 32'd11949, 32'd4924},
{32'd831, 32'd6104, -32'd1032, 32'd6559},
{32'd2825, -32'd2174, -32'd3828, -32'd4457},
{32'd4726, -32'd7483, -32'd3375, 32'd726},
{32'd6273, -32'd558, -32'd1762, -32'd14547},
{-32'd2683, -32'd10196, -32'd3605, -32'd2735},
{-32'd18420, 32'd3153, 32'd1388, 32'd9147},
{-32'd1102, 32'd6503, 32'd4049, 32'd9463},
{32'd12091, 32'd8097, 32'd163, 32'd2665},
{-32'd956, -32'd6239, -32'd1246, -32'd3175}
},
{{32'd4450, 32'd8320, 32'd2436, -32'd3708},
{-32'd13138, -32'd14813, -32'd583, 32'd885},
{-32'd3789, -32'd3801, -32'd1255, -32'd9094},
{32'd7141, 32'd17903, -32'd232, 32'd745},
{32'd800, 32'd9605, 32'd1545, -32'd1490},
{-32'd5657, 32'd4447, -32'd4281, -32'd6339},
{32'd12630, 32'd7047, 32'd829, 32'd2702},
{-32'd89, -32'd244, 32'd1555, 32'd10310},
{32'd448, 32'd7682, 32'd9737, 32'd4322},
{32'd5133, 32'd7098, 32'd5433, 32'd719},
{-32'd885, -32'd10514, -32'd2436, -32'd5705},
{32'd1213, -32'd3936, -32'd8697, 32'd9707},
{-32'd364, 32'd12739, -32'd8505, -32'd3505},
{-32'd751, -32'd6939, 32'd3106, -32'd3933},
{-32'd2839, -32'd5388, -32'd531, 32'd3471},
{-32'd2932, -32'd9880, -32'd3336, -32'd7063},
{32'd4444, 32'd3059, 32'd5258, -32'd1748},
{-32'd10060, -32'd11362, 32'd18489, -32'd146},
{32'd3573, 32'd13606, -32'd12775, -32'd6321},
{-32'd1159, 32'd3346, 32'd1067, -32'd6660},
{32'd9495, -32'd3206, -32'd3676, -32'd8204},
{-32'd2284, -32'd6428, -32'd10266, -32'd7649},
{32'd503, -32'd4883, -32'd2396, 32'd9540},
{-32'd3804, 32'd2691, -32'd3117, 32'd6273},
{32'd4150, 32'd5189, 32'd9541, -32'd2472},
{32'd3035, 32'd19631, -32'd1411, -32'd6136},
{-32'd2973, 32'd788, -32'd5101, 32'd1406},
{32'd11695, 32'd8028, 32'd6028, 32'd812},
{32'd7379, -32'd5866, -32'd4584, -32'd12284},
{32'd4297, -32'd23, -32'd751, -32'd5242},
{-32'd1190, -32'd5817, -32'd6454, -32'd2806},
{32'd2037, -32'd2621, -32'd11152, 32'd1026},
{32'd2582, 32'd9785, 32'd3215, 32'd213},
{-32'd4554, -32'd6323, 32'd2221, 32'd4032},
{32'd3268, 32'd3841, 32'd1060, -32'd5237},
{-32'd926, 32'd150, 32'd755, 32'd1098},
{32'd2908, 32'd2020, 32'd3407, 32'd9148},
{-32'd5015, -32'd2996, 32'd10440, 32'd4091},
{-32'd576, 32'd4435, 32'd6499, 32'd8231},
{-32'd1596, 32'd1173, 32'd7312, 32'd2825},
{-32'd2300, -32'd2286, 32'd2777, 32'd4068},
{-32'd2350, 32'd1997, 32'd4682, -32'd11412},
{-32'd6410, 32'd13675, 32'd5267, -32'd603},
{32'd4516, 32'd526, -32'd10368, 32'd8530},
{-32'd2411, 32'd5390, 32'd7062, -32'd859},
{32'd6155, 32'd748, 32'd5112, 32'd3615},
{32'd4826, -32'd10758, -32'd1668, -32'd5878},
{-32'd12913, -32'd9610, 32'd4913, 32'd13172},
{32'd19038, 32'd1660, -32'd4711, -32'd2053},
{-32'd6378, -32'd3767, 32'd7094, -32'd233},
{32'd1165, 32'd967, 32'd107, -32'd6214},
{32'd8441, -32'd1966, -32'd6701, 32'd6208},
{-32'd7406, -32'd976, -32'd6603, -32'd11961},
{32'd1622, 32'd2861, -32'd7889, -32'd374},
{-32'd1204, 32'd3504, -32'd3602, -32'd880},
{32'd3817, -32'd5676, 32'd3067, 32'd996},
{-32'd3765, -32'd46, 32'd3974, 32'd6912},
{-32'd561, -32'd1289, -32'd5605, -32'd4748},
{-32'd3776, -32'd11182, -32'd1984, 32'd9100},
{-32'd13144, -32'd407, -32'd3049, 32'd1364},
{-32'd6063, 32'd5651, -32'd7081, 32'd4668},
{32'd9208, 32'd2143, 32'd2494, 32'd3268},
{32'd6699, 32'd137, -32'd6732, 32'd310},
{32'd2721, 32'd3685, -32'd1093, -32'd9034},
{32'd1413, -32'd762, 32'd6293, 32'd9300},
{-32'd7592, 32'd11591, -32'd2505, -32'd92},
{-32'd2651, 32'd6046, -32'd2546, 32'd8316},
{32'd5195, 32'd7748, -32'd3096, 32'd3384},
{-32'd3210, -32'd4928, 32'd3755, -32'd954},
{-32'd3467, -32'd3912, -32'd5147, -32'd7288},
{32'd5366, -32'd1623, 32'd258, 32'd1220},
{-32'd5173, -32'd3010, 32'd658, 32'd4466},
{32'd283, -32'd6688, -32'd6064, -32'd4606},
{-32'd3804, -32'd2577, 32'd4243, -32'd6696},
{32'd8167, 32'd6841, 32'd1225, -32'd7595},
{32'd1251, 32'd5613, -32'd1489, 32'd6098},
{-32'd8853, -32'd11110, 32'd10923, -32'd5530},
{32'd15442, -32'd5432, -32'd1490, -32'd2281},
{-32'd1023, 32'd13892, -32'd21, -32'd5838},
{32'd3431, -32'd5778, 32'd3595, 32'd4602},
{32'd1465, 32'd11824, 32'd4852, 32'd5185},
{32'd2925, -32'd2205, 32'd2166, 32'd3},
{-32'd1776, -32'd4266, -32'd9795, -32'd6897},
{-32'd399, -32'd941, 32'd6961, 32'd3124},
{-32'd11579, -32'd2831, -32'd5731, -32'd241},
{-32'd3778, 32'd4424, -32'd7239, 32'd8531},
{-32'd1536, 32'd1135, -32'd197, -32'd8972},
{-32'd2296, -32'd8219, 32'd422, -32'd9775},
{32'd5827, -32'd5101, 32'd3572, 32'd1202},
{-32'd4972, -32'd3379, -32'd2660, -32'd3510},
{-32'd3500, -32'd368, 32'd5813, 32'd1744},
{32'd1182, -32'd2887, -32'd5435, -32'd83},
{-32'd12499, 32'd4279, 32'd4552, 32'd1882},
{-32'd6171, -32'd6880, -32'd1375, -32'd1361},
{32'd2422, -32'd1915, -32'd2287, -32'd13319},
{-32'd2552, -32'd1018, 32'd3271, -32'd3733},
{32'd6179, 32'd3821, 32'd1533, -32'd576},
{-32'd6255, 32'd10580, -32'd418, 32'd13811},
{-32'd807, 32'd668, 32'd929, -32'd9402},
{32'd8874, 32'd8313, 32'd8207, 32'd4643},
{-32'd7561, -32'd2710, -32'd4235, 32'd1081},
{-32'd18806, -32'd12004, -32'd308, -32'd6338},
{32'd7333, 32'd2944, -32'd7585, 32'd6879},
{32'd2367, -32'd8231, 32'd2702, -32'd5544},
{32'd7461, -32'd2234, 32'd4100, 32'd12818},
{32'd2404, -32'd2685, 32'd4735, -32'd9628},
{-32'd1027, -32'd61, 32'd4950, 32'd4324},
{-32'd8834, -32'd4229, -32'd6318, 32'd8966},
{32'd8165, 32'd11193, 32'd926, 32'd1497},
{-32'd7866, -32'd1520, -32'd2667, 32'd7432},
{32'd2572, -32'd3317, -32'd1973, 32'd4137},
{32'd6403, -32'd2979, -32'd6296, -32'd1821},
{-32'd2413, 32'd9257, 32'd5448, -32'd182},
{32'd6071, -32'd3737, -32'd4351, -32'd5593},
{32'd1825, 32'd3904, -32'd6612, -32'd10227},
{-32'd4081, -32'd4019, -32'd3685, -32'd9797},
{-32'd4158, 32'd3219, -32'd6099, 32'd3270},
{-32'd6645, 32'd2755, 32'd4060, 32'd5578},
{-32'd2045, 32'd5930, 32'd14869, 32'd5664},
{32'd5922, 32'd2692, -32'd2765, 32'd4561},
{32'd2693, 32'd10679, -32'd6446, -32'd1838},
{32'd9049, -32'd591, -32'd2329, -32'd1517},
{-32'd7354, -32'd2917, -32'd1062, 32'd14636},
{32'd10, 32'd1676, 32'd7136, -32'd6945},
{32'd571, -32'd1211, -32'd13592, -32'd5342},
{32'd10217, 32'd7747, 32'd3584, -32'd7916},
{-32'd5235, 32'd648, -32'd3561, -32'd3882},
{-32'd5552, -32'd7578, -32'd3776, -32'd6442},
{32'd2144, -32'd5432, -32'd152, -32'd5533},
{32'd3932, -32'd10581, -32'd335, 32'd7685},
{-32'd12408, -32'd3701, -32'd5279, -32'd6655},
{-32'd5124, -32'd7595, 32'd4356, 32'd5475},
{-32'd4008, -32'd2408, -32'd190, -32'd3917},
{32'd3270, 32'd4888, 32'd2539, 32'd8161},
{32'd14877, 32'd12558, 32'd7034, -32'd3693},
{-32'd542, -32'd1871, 32'd222, 32'd431},
{-32'd1651, 32'd6545, 32'd6023, 32'd3490},
{32'd5560, 32'd9062, 32'd3357, 32'd7142},
{-32'd3598, 32'd1496, 32'd1308, -32'd11369},
{-32'd7091, -32'd9205, 32'd4144, 32'd3088},
{32'd10660, 32'd13795, 32'd2398, 32'd548},
{-32'd6152, 32'd2449, 32'd3977, -32'd9540},
{-32'd1065, 32'd3685, -32'd4881, -32'd7160},
{-32'd4235, 32'd4830, -32'd2845, 32'd4039},
{32'd237, 32'd4840, 32'd5041, -32'd6532},
{32'd8185, 32'd2061, 32'd5516, 32'd1886},
{-32'd868, -32'd8839, 32'd853, -32'd1840},
{32'd817, -32'd6933, 32'd8535, 32'd10256},
{-32'd11100, 32'd5414, -32'd986, 32'd4218},
{-32'd13268, -32'd4621, -32'd6154, -32'd11236},
{32'd9054, -32'd3732, 32'd2156, 32'd3848},
{32'd7932, 32'd3717, -32'd6938, 32'd3018},
{-32'd4308, -32'd4324, -32'd9143, -32'd5669},
{-32'd1637, -32'd4128, 32'd7451, -32'd5246},
{-32'd8933, -32'd5298, -32'd1566, 32'd8672},
{-32'd4065, 32'd16684, -32'd2074, -32'd8367},
{32'd2450, -32'd299, 32'd1164, -32'd2485},
{-32'd3058, -32'd6860, 32'd766, 32'd8898},
{-32'd8760, -32'd17583, -32'd4717, -32'd5384},
{32'd121, 32'd6826, 32'd6203, 32'd635},
{32'd6484, 32'd5079, 32'd2670, 32'd561},
{32'd6087, 32'd14289, -32'd1143, 32'd16109},
{32'd7408, -32'd1711, -32'd793, 32'd4181},
{32'd5108, 32'd7548, 32'd4238, -32'd2503},
{-32'd14387, -32'd12418, 32'd4262, 32'd4010},
{-32'd3374, -32'd2083, 32'd574, 32'd1249},
{32'd5140, 32'd8440, 32'd5783, 32'd3978},
{-32'd976, -32'd12154, -32'd81, 32'd3585},
{32'd705, 32'd4406, -32'd1156, -32'd4832},
{-32'd4108, -32'd15858, -32'd5496, -32'd8154},
{-32'd1179, -32'd13706, 32'd12132, -32'd546},
{-32'd616, 32'd156, -32'd1693, -32'd10334},
{32'd3290, 32'd5453, 32'd5338, -32'd9996},
{32'd4060, 32'd5155, 32'd821, -32'd181},
{32'd1681, 32'd6159, -32'd1024, -32'd2652},
{32'd3676, -32'd6927, 32'd2788, 32'd8901},
{32'd3146, -32'd5096, 32'd2622, 32'd7109},
{-32'd5355, 32'd4786, -32'd7167, -32'd2681},
{-32'd702, 32'd1061, -32'd7502, -32'd1864},
{-32'd13887, -32'd1523, -32'd4644, 32'd9024},
{32'd7378, 32'd3311, 32'd1462, 32'd2646},
{32'd2073, -32'd14512, -32'd2213, 32'd9476},
{-32'd3667, -32'd5377, 32'd3246, 32'd2320},
{-32'd2972, -32'd1282, -32'd8227, -32'd7016},
{-32'd6004, -32'd6625, -32'd5479, -32'd1539},
{-32'd1307, -32'd288, 32'd2168, -32'd4232},
{-32'd5284, 32'd7326, -32'd3888, -32'd1138},
{-32'd14653, -32'd5737, 32'd3139, -32'd1724},
{-32'd5258, 32'd3424, 32'd1507, -32'd612},
{32'd30, 32'd1900, 32'd834, 32'd4519},
{-32'd10681, 32'd3297, 32'd289, 32'd6126},
{-32'd5758, -32'd2315, 32'd7718, 32'd5991},
{-32'd8062, -32'd8932, -32'd2462, 32'd548},
{-32'd6754, 32'd6359, 32'd3487, 32'd8675},
{32'd6208, -32'd2465, 32'd7918, -32'd1067},
{32'd3858, 32'd3262, 32'd1503, -32'd3887},
{32'd2705, 32'd824, -32'd104, 32'd9417},
{-32'd5783, -32'd8637, 32'd3570, -32'd526},
{32'd3274, 32'd1376, 32'd1148, 32'd1433},
{-32'd1480, -32'd908, 32'd13584, -32'd1372},
{-32'd2765, -32'd9083, 32'd66, -32'd777},
{-32'd6358, 32'd7011, -32'd8819, 32'd2141},
{32'd53, -32'd6312, -32'd1220, 32'd9559},
{32'd269, 32'd5392, -32'd1080, -32'd10158},
{-32'd1362, -32'd5445, -32'd1745, 32'd1440},
{32'd1363, -32'd1153, 32'd2346, -32'd3866},
{32'd7924, 32'd1374, 32'd1361, -32'd4920},
{32'd770, -32'd5447, 32'd2138, -32'd2875},
{32'd15224, -32'd4128, 32'd3830, -32'd2067},
{32'd2670, 32'd4681, 32'd2456, 32'd460},
{-32'd3231, -32'd12790, -32'd1856, 32'd9607},
{32'd7075, -32'd9719, 32'd4075, 32'd7242},
{-32'd4152, 32'd4589, -32'd1318, -32'd2776},
{-32'd2439, -32'd4377, 32'd4380, 32'd460},
{32'd6069, 32'd920, -32'd1591, 32'd4535},
{-32'd14530, -32'd4612, -32'd8734, -32'd1128},
{-32'd5268, -32'd1367, 32'd3016, -32'd6454},
{-32'd1166, 32'd4968, -32'd8265, 32'd9558},
{32'd162, -32'd4473, 32'd10847, -32'd2442},
{32'd542, 32'd6311, 32'd4396, 32'd6580},
{32'd4118, -32'd3795, 32'd9686, 32'd9873},
{32'd2806, 32'd3025, -32'd9329, -32'd87},
{32'd8180, 32'd3133, -32'd4069, -32'd2734},
{-32'd6937, -32'd12521, -32'd17228, -32'd3873},
{32'd181, 32'd6579, -32'd11813, -32'd3736},
{-32'd6654, -32'd2344, 32'd8806, -32'd19245},
{32'd4805, -32'd5730, 32'd1644, -32'd2430},
{-32'd22920, 32'd1183, 32'd911, -32'd1954},
{-32'd1477, 32'd3113, -32'd146, -32'd8776},
{32'd4940, 32'd17950, 32'd6139, 32'd8470},
{-32'd1119, -32'd14912, -32'd2217, -32'd7893},
{32'd3077, 32'd3400, -32'd9206, 32'd1836},
{-32'd1819, -32'd7361, 32'd2121, -32'd5926},
{32'd8787, 32'd9416, -32'd6313, 32'd3112},
{32'd3559, 32'd2335, 32'd1367, 32'd5995},
{-32'd5035, 32'd8179, -32'd2328, 32'd4068},
{-32'd3971, -32'd8363, 32'd3146, -32'd1223},
{32'd8493, 32'd906, -32'd5190, 32'd5310},
{32'd1377, 32'd14945, 32'd455, 32'd4287},
{32'd844, -32'd4880, 32'd4651, 32'd1482},
{-32'd3975, 32'd8275, -32'd6516, -32'd9788},
{32'd3912, 32'd7244, 32'd3008, -32'd5828},
{32'd2370, 32'd1851, -32'd912, 32'd1520},
{-32'd5768, 32'd72, 32'd10587, 32'd2388},
{32'd10850, 32'd7258, 32'd3253, -32'd4901},
{32'd3136, -32'd526, -32'd3200, -32'd7929},
{-32'd5761, -32'd3917, 32'd6168, 32'd5317},
{-32'd1253, -32'd7348, 32'd3486, 32'd1408},
{32'd589, -32'd6889, 32'd3502, -32'd4996},
{32'd3058, -32'd7269, 32'd2535, -32'd7090},
{-32'd8659, -32'd10245, 32'd7407, 32'd2584},
{32'd5933, 32'd742, -32'd3519, 32'd4793},
{32'd7886, 32'd12044, 32'd1199, 32'd2132},
{32'd6311, 32'd1075, -32'd3380, -32'd9945},
{-32'd1837, -32'd2505, -32'd4967, 32'd293},
{-32'd2079, -32'd4481, 32'd2076, -32'd13707},
{32'd7118, -32'd3819, 32'd660, 32'd2298},
{32'd1762, 32'd9840, -32'd647, -32'd1355},
{-32'd6355, -32'd10453, -32'd6907, -32'd3262},
{32'd9209, 32'd3858, 32'd10784, 32'd2164},
{-32'd5767, -32'd7173, -32'd1351, -32'd5357},
{32'd8039, 32'd4718, -32'd3998, 32'd2645},
{32'd658, 32'd3355, -32'd739, -32'd202},
{32'd12337, -32'd243, 32'd9580, -32'd4615},
{-32'd7785, -32'd1514, 32'd2177, 32'd11123},
{-32'd2329, -32'd5978, -32'd1991, -32'd4186},
{-32'd2339, 32'd8422, -32'd4411, 32'd3218},
{-32'd10861, 32'd2881, 32'd4095, 32'd11027},
{-32'd14324, -32'd10699, -32'd2720, 32'd2825},
{32'd4119, -32'd8473, -32'd6528, -32'd1503},
{32'd2298, -32'd3424, 32'd1622, 32'd163},
{32'd737, 32'd5242, -32'd5747, 32'd2659},
{32'd10079, -32'd5198, -32'd5347, 32'd4414},
{-32'd4069, 32'd1756, -32'd3019, 32'd8080},
{-32'd6647, -32'd2121, 32'd7069, -32'd5439},
{32'd2276, -32'd6042, -32'd1462, 32'd5775},
{32'd3899, 32'd7009, 32'd3842, 32'd339},
{32'd2010, -32'd243, 32'd2635, -32'd3186},
{-32'd6403, -32'd3848, 32'd1698, 32'd3404},
{-32'd1547, 32'd4471, 32'd1991, 32'd12058},
{32'd2079, 32'd8247, -32'd1637, 32'd10847},
{32'd3584, -32'd5786, 32'd10269, 32'd1992},
{32'd8052, 32'd484, 32'd4909, -32'd3922},
{32'd9201, 32'd1960, 32'd7410, -32'd3284},
{-32'd1563, -32'd7161, 32'd2202, -32'd1760},
{32'd1723, -32'd3441, -32'd4710, 32'd6735},
{32'd2052, 32'd7791, -32'd5444, 32'd2601},
{32'd6522, -32'd4023, -32'd1729, 32'd19570},
{32'd5706, 32'd4223, 32'd17710, 32'd4986},
{32'd2921, -32'd1430, -32'd3180, 32'd8470},
{-32'd6168, -32'd6241, -32'd3361, -32'd1256},
{32'd1662, 32'd1988, 32'd1749, -32'd1575},
{32'd130, -32'd9770, -32'd1773, 32'd1845},
{32'd137, -32'd6463, -32'd743, 32'd8019},
{-32'd6774, 32'd916, -32'd6166, 32'd11254},
{32'd816, -32'd1926, 32'd1247, 32'd3646},
{-32'd6199, -32'd3938, 32'd6083, -32'd6972},
{-32'd7406, -32'd458, -32'd10043, -32'd5068},
{-32'd25, 32'd3671, 32'd2083, -32'd3067},
{32'd6550, -32'd1725, -32'd4531, -32'd5946}
},
{{-32'd3085, -32'd4126, -32'd7478, -32'd1731},
{-32'd11739, -32'd10550, -32'd943, -32'd3889},
{-32'd5489, 32'd6459, 32'd10383, -32'd14021},
{32'd7726, 32'd6876, -32'd4560, -32'd2631},
{32'd3277, 32'd3821, 32'd5717, -32'd4234},
{-32'd1641, 32'd7345, -32'd7626, -32'd4478},
{32'd2355, 32'd539, 32'd3160, 32'd10363},
{-32'd1531, 32'd3710, -32'd8996, -32'd5312},
{32'd8911, -32'd7199, 32'd4395, -32'd9110},
{32'd4947, 32'd7434, -32'd3178, -32'd1777},
{32'd5662, -32'd735, 32'd7598, -32'd7182},
{32'd8857, 32'd2926, -32'd8750, -32'd11945},
{-32'd6449, 32'd7597, 32'd837, 32'd4074},
{-32'd8719, -32'd7699, -32'd11963, -32'd4913},
{-32'd7237, -32'd676, -32'd12098, -32'd17312},
{32'd3264, -32'd492, -32'd4481, -32'd4971},
{-32'd3699, -32'd2564, 32'd5858, 32'd4052},
{-32'd5002, 32'd4261, -32'd7493, -32'd6951},
{32'd5964, 32'd4558, 32'd2389, -32'd2509},
{32'd2652, -32'd11860, 32'd13386, 32'd378},
{-32'd3044, -32'd2757, 32'd2508, -32'd5935},
{-32'd3656, -32'd10054, 32'd2720, -32'd6977},
{-32'd14352, -32'd12766, -32'd17243, 32'd9106},
{32'd2676, 32'd6374, -32'd5576, 32'd2689},
{32'd6975, 32'd13326, -32'd8558, 32'd5234},
{32'd6553, 32'd9680, -32'd1520, -32'd7628},
{-32'd4701, -32'd2573, -32'd5964, 32'd5243},
{-32'd6480, 32'd2207, 32'd9139, 32'd1911},
{32'd6114, 32'd1251, -32'd8123, 32'd10106},
{32'd647, 32'd1151, 32'd3164, 32'd10438},
{-32'd9970, 32'd5934, -32'd5593, -32'd8948},
{32'd2131, -32'd7004, 32'd3689, 32'd16753},
{32'd6886, 32'd11304, 32'd1970, 32'd17311},
{32'd33, 32'd9235, -32'd3681, -32'd10319},
{-32'd670, 32'd1646, 32'd433, -32'd4351},
{32'd10313, 32'd7260, 32'd3292, -32'd12408},
{-32'd12758, -32'd4061, 32'd3033, 32'd6977},
{32'd12711, 32'd11070, -32'd3468, -32'd1416},
{32'd972, -32'd2662, 32'd4047, 32'd7969},
{-32'd2834, -32'd5021, 32'd8988, 32'd6035},
{32'd15474, -32'd4329, 32'd3314, -32'd1237},
{32'd4768, -32'd3647, 32'd10646, 32'd2985},
{-32'd3663, -32'd7852, 32'd10172, -32'd4352},
{-32'd9984, 32'd170, -32'd13736, -32'd8713},
{-32'd6501, -32'd5226, -32'd4522, -32'd6452},
{-32'd6682, -32'd4377, 32'd942, -32'd6338},
{32'd5277, -32'd2102, -32'd4728, -32'd8564},
{-32'd3074, 32'd4972, -32'd3823, -32'd358},
{-32'd7537, 32'd4820, -32'd11320, -32'd8367},
{-32'd11901, -32'd12663, 32'd1261, 32'd12218},
{-32'd12989, -32'd12755, 32'd891, 32'd983},
{-32'd3776, 32'd10438, -32'd8794, -32'd2020},
{32'd2020, -32'd12994, -32'd11876, -32'd12887},
{32'd154, 32'd3064, 32'd11953, 32'd16259},
{32'd1683, 32'd6386, -32'd17913, 32'd1250},
{-32'd14052, -32'd8845, 32'd1278, -32'd3001},
{32'd1484, 32'd64, 32'd7297, 32'd11557},
{-32'd4956, -32'd4205, 32'd3337, 32'd6373},
{32'd5931, -32'd4313, -32'd9627, -32'd12002},
{-32'd10426, -32'd19657, -32'd5953, 32'd4745},
{32'd2072, 32'd4704, -32'd8319, -32'd361},
{32'd17583, -32'd3540, 32'd2093, 32'd6375},
{-32'd3446, -32'd10472, 32'd17921, 32'd2039},
{-32'd3011, -32'd12461, 32'd775, 32'd4250},
{32'd386, -32'd896, -32'd119, -32'd3158},
{-32'd1989, -32'd618, 32'd1521, -32'd10402},
{-32'd9754, 32'd4790, -32'd10230, -32'd12592},
{-32'd7684, -32'd10538, -32'd16937, -32'd17361},
{32'd13796, 32'd6112, 32'd4262, -32'd6849},
{-32'd4263, -32'd2338, -32'd5911, -32'd154},
{-32'd4361, -32'd12245, -32'd1914, -32'd5444},
{-32'd10845, 32'd1101, -32'd13561, -32'd8692},
{-32'd5833, 32'd3168, 32'd9286, 32'd582},
{-32'd4471, 32'd2344, 32'd3643, 32'd8316},
{32'd11461, 32'd6606, 32'd4499, 32'd5472},
{-32'd5711, 32'd6499, 32'd3611, 32'd8673},
{-32'd15630, 32'd6934, 32'd1894, 32'd701},
{-32'd1703, -32'd735, 32'd3081, 32'd3399},
{-32'd3682, 32'd2939, 32'd149, 32'd5004},
{-32'd9953, 32'd1137, -32'd6256, 32'd4448},
{32'd17209, 32'd7938, 32'd234, 32'd5942},
{32'd1044, -32'd334, 32'd14086, -32'd2636},
{-32'd11543, 32'd5298, 32'd15530, 32'd6741},
{-32'd13519, 32'd632, 32'd1192, 32'd3215},
{32'd2093, -32'd9010, -32'd15154, 32'd3140},
{-32'd4284, -32'd16705, 32'd8993, -32'd16241},
{32'd5169, 32'd4379, 32'd5941, -32'd4372},
{-32'd5798, -32'd3509, 32'd5970, 32'd5603},
{32'd7723, -32'd12545, 32'd14323, -32'd4185},
{-32'd12001, -32'd10337, 32'd3869, -32'd12556},
{32'd5181, 32'd2679, -32'd1303, -32'd1403},
{-32'd1969, -32'd11732, 32'd6011, 32'd2638},
{32'd5116, 32'd5410, -32'd19096, -32'd13031},
{-32'd2281, -32'd5392, 32'd2783, -32'd3304},
{32'd3581, 32'd4350, -32'd2496, -32'd8646},
{-32'd5685, 32'd1647, -32'd1504, -32'd7669},
{32'd25279, 32'd5924, 32'd1594, -32'd1669},
{32'd421, 32'd8744, -32'd5060, 32'd717},
{32'd10164, 32'd169, 32'd14272, 32'd10097},
{32'd4710, 32'd8755, -32'd273, -32'd8173},
{-32'd8272, -32'd9304, -32'd15566, -32'd18766},
{-32'd10084, -32'd12332, 32'd716, 32'd3610},
{32'd10863, 32'd5752, -32'd3134, 32'd9265},
{32'd235, 32'd10190, -32'd6401, 32'd2777},
{-32'd4992, -32'd2996, 32'd698, 32'd4659},
{32'd1172, 32'd3037, -32'd12598, -32'd12158},
{32'd3067, 32'd1073, 32'd655, 32'd7621},
{-32'd5056, -32'd7187, 32'd5131, 32'd10361},
{-32'd5571, 32'd11189, -32'd2102, -32'd5987},
{-32'd6945, -32'd10531, 32'd14472, -32'd2514},
{32'd939, -32'd8568, 32'd5174, -32'd2147},
{32'd12906, -32'd4331, 32'd15459, 32'd4851},
{32'd7425, 32'd4627, 32'd25472, 32'd11968},
{32'd14312, 32'd11884, 32'd4578, -32'd1427},
{32'd5242, -32'd8894, -32'd4316, -32'd1089},
{32'd1161, -32'd12136, -32'd8007, 32'd9674},
{-32'd1521, -32'd4050, -32'd10762, -32'd3447},
{32'd8359, 32'd11654, -32'd3338, 32'd13045},
{32'd1140, 32'd5667, 32'd583, 32'd2665},
{-32'd2442, -32'd1600, -32'd6227, -32'd12872},
{-32'd11806, 32'd1231, -32'd1561, -32'd11888},
{32'd11982, 32'd2696, 32'd7863, -32'd10602},
{-32'd10709, 32'd5867, -32'd10522, -32'd9486},
{32'd4177, 32'd2880, -32'd973, -32'd2287},
{32'd3617, 32'd2448, 32'd4888, 32'd9385},
{-32'd9910, 32'd5104, -32'd4795, 32'd4914},
{32'd5569, -32'd6611, -32'd3072, -32'd5015},
{-32'd948, -32'd9632, -32'd2033, -32'd13408},
{32'd4044, 32'd5039, -32'd3469, -32'd8869},
{32'd222, -32'd7668, -32'd8297, 32'd8696},
{32'd5186, 32'd18891, 32'd12412, 32'd3228},
{32'd3762, -32'd381, -32'd7302, 32'd13558},
{-32'd6483, -32'd870, 32'd96, 32'd429},
{-32'd1795, 32'd6915, -32'd10756, 32'd10052},
{32'd13152, 32'd459, 32'd175, -32'd327},
{32'd5465, -32'd8450, 32'd9966, 32'd10976},
{-32'd7337, 32'd187, -32'd4296, 32'd3140},
{-32'd1204, -32'd6936, 32'd1116, -32'd7471},
{32'd9490, 32'd7754, 32'd3348, 32'd5990},
{-32'd8063, -32'd17619, -32'd10800, 32'd1924},
{-32'd6974, -32'd987, 32'd3858, 32'd8880},
{-32'd56, -32'd3450, -32'd6586, -32'd8056},
{-32'd8759, -32'd7896, -32'd3520, -32'd3505},
{32'd2787, -32'd6663, -32'd15596, 32'd8171},
{32'd1908, 32'd3102, -32'd4530, -32'd5730},
{-32'd12970, -32'd739, -32'd117, 32'd2277},
{-32'd3440, -32'd21257, 32'd10418, -32'd12276},
{-32'd3711, -32'd8394, 32'd11382, 32'd7826},
{32'd14515, -32'd845, -32'd163, 32'd20256},
{-32'd12367, 32'd6071, -32'd566, 32'd7979},
{-32'd1685, 32'd3970, -32'd1445, 32'd337},
{32'd173, 32'd7875, -32'd7207, 32'd7746},
{-32'd580, -32'd2701, 32'd1605, -32'd3210},
{-32'd8011, -32'd1531, 32'd1221, -32'd1842},
{-32'd4146, -32'd7927, 32'd5124, 32'd11987},
{32'd8315, -32'd733, -32'd6736, -32'd614},
{32'd6521, 32'd1975, 32'd8316, 32'd21},
{-32'd13128, 32'd8537, -32'd13332, 32'd1653},
{32'd2849, -32'd2850, 32'd1122, 32'd2759},
{32'd1152, -32'd2337, 32'd7670, -32'd7970},
{-32'd317, 32'd9883, 32'd11607, -32'd11282},
{-32'd5526, 32'd4076, -32'd14419, -32'd17418},
{32'd13960, -32'd11378, 32'd5777, -32'd1672},
{32'd9169, 32'd11077, 32'd15060, -32'd3166},
{-32'd5014, -32'd980, 32'd5740, -32'd8619},
{-32'd834, 32'd1335, 32'd6977, 32'd23176},
{-32'd11017, 32'd3756, -32'd22215, 32'd4574},
{32'd9809, -32'd5521, -32'd3578, -32'd18},
{-32'd1205, -32'd5737, 32'd13572, 32'd5277},
{32'd1213, -32'd466, -32'd6592, 32'd5255},
{32'd3549, 32'd5679, -32'd2907, 32'd17997},
{-32'd10676, 32'd9411, -32'd11745, 32'd18739},
{32'd5627, 32'd4182, -32'd710, 32'd3679},
{-32'd2472, 32'd5243, -32'd13344, -32'd4073},
{32'd10619, -32'd323, 32'd894, 32'd11662},
{-32'd1407, 32'd6021, 32'd2694, -32'd16381},
{-32'd2333, 32'd8786, 32'd9539, 32'd5908},
{-32'd512, -32'd564, -32'd1141, -32'd2203},
{32'd10328, 32'd622, -32'd8881, 32'd5820},
{-32'd7722, 32'd346, 32'd2764, -32'd3391},
{32'd3048, 32'd915, -32'd10439, 32'd1481},
{-32'd5801, -32'd11254, 32'd6425, 32'd5226},
{-32'd14799, -32'd2928, -32'd2284, 32'd2031},
{-32'd2304, -32'd6418, 32'd12177, 32'd101},
{-32'd17237, -32'd3816, -32'd17880, -32'd4970},
{32'd3353, 32'd3282, -32'd5608, -32'd6397},
{32'd5771, 32'd3672, -32'd1549, 32'd2709},
{32'd13481, -32'd3291, -32'd2098, 32'd2824},
{-32'd14549, -32'd3884, 32'd6785, 32'd19507},
{-32'd725, 32'd210, -32'd11504, 32'd539},
{32'd2205, 32'd4112, -32'd1779, 32'd9404},
{32'd2322, -32'd1145, 32'd1394, 32'd7971},
{-32'd12716, -32'd5195, 32'd824, -32'd6825},
{-32'd8277, -32'd11307, -32'd4339, 32'd13268},
{32'd2773, -32'd16115, -32'd2802, -32'd16143},
{-32'd6941, -32'd7571, -32'd23795, 32'd2019},
{-32'd5542, -32'd6318, -32'd11428, 32'd8131},
{-32'd4740, -32'd3976, -32'd3778, 32'd1096},
{-32'd3053, 32'd3194, -32'd2841, -32'd532},
{-32'd8720, -32'd469, -32'd2705, -32'd12718},
{-32'd3590, -32'd6234, 32'd1605, -32'd5790},
{32'd1144, 32'd8687, 32'd3201, 32'd2878},
{32'd2439, -32'd2674, 32'd23944, 32'd10119},
{32'd3417, 32'd13831, 32'd10675, 32'd8562},
{-32'd3332, 32'd2752, 32'd15529, -32'd22176},
{32'd1020, 32'd2371, -32'd15198, 32'd8646},
{32'd670, 32'd3954, 32'd2570, -32'd9784},
{-32'd6676, -32'd274, -32'd5218, 32'd2316},
{32'd546, 32'd1378, 32'd5881, -32'd2962},
{32'd2042, -32'd2132, 32'd4437, -32'd13987},
{-32'd9729, -32'd12456, -32'd3106, -32'd13933},
{-32'd7328, -32'd8589, -32'd4112, -32'd8012},
{-32'd3378, -32'd2291, 32'd1492, 32'd157},
{32'd15270, 32'd1258, -32'd8849, -32'd6487},
{-32'd7232, -32'd19375, 32'd11381, -32'd5239},
{-32'd6601, -32'd7693, -32'd18500, 32'd10014},
{32'd3121, -32'd13663, 32'd6549, -32'd7136},
{-32'd3989, 32'd13687, -32'd9486, 32'd13410},
{32'd5258, 32'd6004, 32'd6107, 32'd15181},
{32'd15178, 32'd1068, -32'd443, -32'd2788},
{32'd3435, -32'd6666, 32'd1904, -32'd7777},
{32'd3221, 32'd817, -32'd865, 32'd5326},
{32'd7079, -32'd1067, -32'd3126, -32'd2234},
{32'd10751, -32'd8297, -32'd6464, 32'd6880},
{-32'd8460, -32'd449, 32'd6899, -32'd7610},
{-32'd2338, -32'd4245, 32'd3856, -32'd2348},
{32'd11327, 32'd6473, -32'd2213, -32'd3613},
{-32'd15097, -32'd17004, 32'd1965, -32'd4099},
{32'd6354, 32'd5612, 32'd3258, 32'd5226},
{-32'd12625, 32'd4690, 32'd12056, -32'd2428},
{32'd2224, -32'd1411, 32'd7524, -32'd5780},
{32'd3456, -32'd4166, -32'd17077, -32'd5070},
{32'd2089, -32'd2147, 32'd7640, -32'd4611},
{-32'd16495, -32'd8537, -32'd7240, -32'd12441},
{-32'd6515, 32'd4231, 32'd1515, 32'd1013},
{32'd267, 32'd1878, -32'd9187, -32'd12634},
{32'd8251, 32'd5670, -32'd9615, -32'd9076},
{-32'd7528, -32'd2003, -32'd12293, 32'd1005},
{32'd6017, 32'd6241, -32'd1343, -32'd638},
{32'd6318, 32'd6297, 32'd8358, -32'd2835},
{32'd1054, -32'd7368, -32'd395, -32'd4934},
{32'd8318, -32'd7938, -32'd7254, -32'd11543},
{-32'd15448, 32'd1685, -32'd1895, 32'd2094},
{-32'd12647, -32'd9303, 32'd10078, -32'd3491},
{32'd1390, 32'd8090, 32'd12311, -32'd5609},
{-32'd2643, 32'd4558, -32'd11570, -32'd731},
{-32'd3323, 32'd2696, 32'd6007, 32'd14842},
{-32'd14354, 32'd5623, -32'd9559, -32'd1421},
{32'd5030, 32'd9700, -32'd8792, -32'd16372},
{-32'd1350, 32'd1874, 32'd2934, -32'd365},
{-32'd4656, 32'd205, 32'd6348, -32'd4792},
{32'd5331, -32'd1963, -32'd12786, 32'd5421},
{32'd8727, 32'd4020, -32'd3608, 32'd5485},
{-32'd5042, 32'd50, 32'd7109, -32'd9458},
{32'd4474, 32'd3813, 32'd15890, 32'd14025},
{32'd1482, -32'd3748, 32'd1858, 32'd7800},
{32'd1966, 32'd7182, -32'd8353, 32'd3330},
{-32'd136, 32'd150, 32'd6427, -32'd1957},
{32'd5348, -32'd1273, 32'd3448, 32'd2980},
{32'd3149, 32'd10294, -32'd2486, -32'd280},
{-32'd653, -32'd2505, -32'd10710, 32'd2801},
{32'd12602, 32'd14358, 32'd4293, -32'd11777},
{32'd6908, -32'd9451, -32'd4684, -32'd3616},
{32'd8600, 32'd5850, -32'd6045, 32'd9560},
{-32'd12419, -32'd4661, -32'd371, -32'd6370},
{32'd8552, -32'd3712, 32'd9293, 32'd5721},
{-32'd2128, 32'd11303, -32'd870, 32'd4433},
{-32'd20056, -32'd8170, 32'd11512, -32'd7030},
{32'd4631, -32'd10398, -32'd5152, -32'd8599},
{-32'd4882, 32'd1537, 32'd8110, 32'd7919},
{32'd3694, 32'd5222, -32'd3003, 32'd379},
{-32'd8922, 32'd5260, -32'd5528, -32'd108},
{32'd7023, -32'd2249, 32'd1427, 32'd2219},
{-32'd7304, -32'd14619, -32'd356, -32'd1897},
{-32'd2632, 32'd8819, -32'd1114, -32'd10155},
{32'd4915, -32'd14999, -32'd2864, 32'd3304},
{32'd6217, 32'd4735, -32'd1530, -32'd2614},
{32'd8200, 32'd16428, -32'd6139, -32'd1919},
{32'd490, -32'd385, 32'd4024, 32'd1015},
{-32'd5700, 32'd7116, -32'd4282, 32'd363},
{32'd1631, -32'd4639, -32'd1792, -32'd5810},
{32'd8512, -32'd10013, 32'd9160, 32'd4923},
{32'd10210, -32'd1909, -32'd2271, 32'd488},
{-32'd7813, 32'd3119, 32'd6120, 32'd7599},
{32'd4518, -32'd8807, 32'd6682, 32'd1981},
{-32'd1965, -32'd7839, 32'd13098, 32'd13753},
{-32'd14559, -32'd937, -32'd926, 32'd1225},
{32'd2040, -32'd13140, 32'd108, -32'd6602},
{32'd3345, 32'd1148, -32'd1419, -32'd7821},
{-32'd1790, -32'd9004, -32'd2552, 32'd4953},
{-32'd4990, -32'd3750, -32'd14317, -32'd6901},
{32'd5120, 32'd1146, 32'd10681, 32'd10052},
{-32'd10408, -32'd7861, -32'd5557, -32'd2970},
{-32'd601, -32'd10419, -32'd1439, -32'd3553},
{32'd12333, -32'd5965, 32'd1602, 32'd7754},
{32'd2667, 32'd6771, -32'd2945, 32'd940},
{-32'd10951, -32'd2269, -32'd16001, -32'd1157},
{32'd15190, -32'd4769, 32'd3347, -32'd3818},
{32'd9669, 32'd905, -32'd5756, 32'd2556},
{-32'd399, 32'd805, 32'd5730, 32'd3143}
},
{{32'd10755, 32'd6610, -32'd1302, 32'd898},
{-32'd17785, 32'd5622, -32'd3024, -32'd5281},
{32'd10957, 32'd7570, -32'd6055, 32'd12710},
{32'd3203, 32'd88, -32'd334, -32'd10127},
{32'd18307, 32'd13821, -32'd9597, -32'd9974},
{-32'd8150, 32'd5167, -32'd3459, 32'd10379},
{32'd1642, -32'd9744, 32'd9064, -32'd4593},
{32'd4913, 32'd5816, 32'd363, 32'd1734},
{32'd100, -32'd9303, 32'd5324, 32'd7053},
{32'd5924, -32'd907, 32'd2050, 32'd3695},
{-32'd2258, 32'd2611, -32'd2264, -32'd1321},
{32'd4829, 32'd14969, 32'd12888, 32'd1948},
{32'd2917, -32'd2554, -32'd1140, -32'd9119},
{-32'd9162, 32'd2327, 32'd3877, -32'd141},
{32'd224, 32'd7371, -32'd8484, 32'd5760},
{-32'd7343, -32'd13157, -32'd1264, -32'd10839},
{32'd11068, 32'd1033, 32'd4975, -32'd4511},
{32'd4809, -32'd6743, 32'd2033, 32'd1299},
{-32'd19530, 32'd14874, -32'd1002, 32'd14127},
{-32'd982, 32'd2445, -32'd3031, 32'd11420},
{-32'd4879, 32'd102, -32'd634, 32'd3555},
{-32'd13568, 32'd3078, 32'd349, 32'd11596},
{32'd7775, 32'd5537, -32'd17909, 32'd4803},
{-32'd3322, 32'd9669, -32'd2834, 32'd2992},
{32'd5733, -32'd1111, -32'd7020, 32'd2976},
{-32'd6750, -32'd3039, -32'd3160, 32'd282},
{-32'd345, 32'd8588, -32'd1263, 32'd10330},
{-32'd2705, -32'd10674, 32'd3250, 32'd5934},
{-32'd2168, 32'd5438, 32'd8513, 32'd2277},
{-32'd2494, 32'd12785, 32'd1785, 32'd1231},
{-32'd5215, 32'd856, -32'd10793, 32'd5441},
{32'd5193, -32'd3902, 32'd17676, 32'd3693},
{-32'd1765, 32'd464, 32'd11860, -32'd1434},
{-32'd8939, -32'd1782, 32'd5069, -32'd10568},
{32'd1960, 32'd7041, -32'd2108, 32'd1315},
{-32'd462, -32'd11397, -32'd11971, -32'd4429},
{32'd2310, -32'd12323, 32'd1496, 32'd1708},
{-32'd5288, -32'd4870, 32'd9106, -32'd20507},
{32'd2110, 32'd6252, -32'd2739, 32'd676},
{32'd2400, 32'd13693, 32'd13581, -32'd4448},
{32'd3118, 32'd2282, 32'd1774, -32'd4128},
{32'd13, -32'd11372, -32'd1600, 32'd1887},
{32'd12275, 32'd2730, 32'd2663, -32'd4860},
{32'd2339, 32'd1918, -32'd4197, -32'd8832},
{-32'd6618, 32'd10373, -32'd8631, 32'd6055},
{-32'd7642, -32'd4419, -32'd665, -32'd13232},
{-32'd13011, -32'd2462, 32'd9468, 32'd9184},
{-32'd3962, -32'd81, 32'd352, 32'd2555},
{-32'd238, 32'd5869, -32'd6539, 32'd4464},
{-32'd5774, 32'd2289, 32'd10803, -32'd8555},
{32'd3699, 32'd4672, 32'd5646, 32'd11820},
{-32'd5321, -32'd4267, 32'd32, -32'd5056},
{32'd8964, 32'd4158, 32'd6273, 32'd3196},
{32'd9029, 32'd20294, -32'd1418, -32'd8738},
{32'd18248, 32'd12978, -32'd8214, -32'd6467},
{-32'd11579, -32'd5476, -32'd2758, 32'd6677},
{32'd5260, 32'd9800, 32'd12950, -32'd6714},
{32'd943, 32'd13866, -32'd15049, 32'd2527},
{32'd1547, 32'd2072, 32'd2844, -32'd1971},
{-32'd1527, -32'd6769, -32'd1051, 32'd58},
{-32'd3475, 32'd1785, -32'd17552, 32'd1836},
{-32'd9508, -32'd6326, 32'd5236, -32'd5758},
{-32'd14469, 32'd5424, -32'd376, 32'd15812},
{32'd42, -32'd9882, -32'd2902, 32'd1677},
{-32'd5384, 32'd13211, -32'd4064, -32'd4227},
{32'd8617, 32'd3458, 32'd923, 32'd3041},
{-32'd2498, -32'd4723, 32'd5618, 32'd551},
{32'd8720, 32'd2065, -32'd1224, -32'd433},
{-32'd5026, 32'd8717, -32'd2625, 32'd1465},
{-32'd3607, 32'd4724, 32'd1429, 32'd10838},
{32'd9384, 32'd4417, -32'd4183, -32'd2891},
{-32'd9412, -32'd10202, 32'd5630, -32'd890},
{-32'd19965, -32'd4204, 32'd8422, 32'd387},
{-32'd794, 32'd527, 32'd6483, -32'd16060},
{32'd8908, 32'd8184, -32'd1526, -32'd3379},
{32'd618, 32'd10419, 32'd11641, -32'd2217},
{-32'd10559, 32'd3143, -32'd14310, -32'd49},
{-32'd2826, 32'd2383, -32'd1302, 32'd1739},
{32'd769, -32'd8136, 32'd8880, 32'd760},
{32'd12223, -32'd11492, -32'd943, -32'd6759},
{32'd9676, -32'd5927, -32'd4833, -32'd7964},
{32'd3672, -32'd8151, -32'd1193, -32'd13135},
{-32'd12397, -32'd813, 32'd866, 32'd3626},
{32'd12464, -32'd7155, -32'd299, -32'd4088},
{32'd2798, 32'd3163, 32'd2990, -32'd12939},
{32'd6513, -32'd10075, -32'd7265, 32'd2313},
{32'd6226, 32'd14665, 32'd3183, 32'd5325},
{-32'd12156, 32'd2552, -32'd8358, 32'd16073},
{-32'd5244, 32'd19411, -32'd19222, -32'd2612},
{-32'd454, 32'd6657, 32'd5336, -32'd2711},
{-32'd2863, 32'd4540, 32'd9351, -32'd1064},
{-32'd8112, -32'd1214, -32'd4002, 32'd94},
{-32'd10451, 32'd3007, -32'd10024, 32'd1557},
{32'd16021, -32'd3624, 32'd3512, -32'd7438},
{32'd4988, -32'd13556, 32'd6686, -32'd1915},
{32'd2722, 32'd21546, -32'd9594, 32'd7342},
{32'd7447, 32'd2391, -32'd2676, -32'd968},
{32'd5028, -32'd10640, -32'd8987, 32'd11757},
{32'd5786, -32'd11372, -32'd2361, -32'd3204},
{32'd16317, -32'd1918, -32'd2737, 32'd159},
{32'd3750, -32'd8360, -32'd11396, 32'd2766},
{-32'd8404, -32'd11929, -32'd7431, 32'd6762},
{32'd7852, 32'd9524, 32'd5208, 32'd5601},
{-32'd4159, 32'd9903, -32'd1198, -32'd7101},
{-32'd4538, -32'd19532, -32'd2031, -32'd9829},
{32'd16301, -32'd2984, -32'd14541, 32'd6776},
{32'd2758, -32'd22658, -32'd8368, -32'd4866},
{32'd1344, -32'd2205, 32'd1663, -32'd13779},
{32'd11945, 32'd5688, -32'd5256, -32'd4962},
{32'd6810, -32'd3147, 32'd808, 32'd2455},
{32'd704, 32'd13207, -32'd5656, -32'd1352},
{-32'd664, 32'd8527, 32'd1684, -32'd1889},
{-32'd1267, 32'd7752, 32'd11903, -32'd8226},
{-32'd2707, 32'd4937, 32'd8460, -32'd1900},
{32'd9454, -32'd13510, -32'd20210, 32'd3553},
{-32'd1052, -32'd6555, 32'd2963, 32'd12605},
{32'd5332, -32'd1478, -32'd3228, 32'd4179},
{32'd994, 32'd1764, -32'd4899, -32'd3210},
{32'd2665, -32'd16512, 32'd10248, -32'd5935},
{-32'd2413, -32'd11803, 32'd10053, 32'd9826},
{32'd5330, 32'd5294, -32'd2307, 32'd1658},
{-32'd11210, 32'd6704, -32'd1928, -32'd2354},
{-32'd2358, -32'd901, 32'd1409, -32'd16309},
{32'd3844, 32'd7476, -32'd10999, 32'd6441},
{-32'd2144, 32'd20100, -32'd1202, 32'd1843},
{32'd3476, 32'd11546, 32'd8203, 32'd11339},
{32'd568, -32'd18276, -32'd2208, 32'd3827},
{-32'd5182, 32'd4831, -32'd9849, 32'd3665},
{32'd7419, -32'd9819, -32'd2490, 32'd5181},
{-32'd2086, 32'd13675, 32'd3466, -32'd8664},
{32'd4965, -32'd9541, 32'd4428, -32'd6107},
{32'd1652, 32'd6317, 32'd8960, 32'd1666},
{-32'd6886, 32'd733, -32'd1073, 32'd550},
{32'd3445, -32'd11889, 32'd5344, 32'd2272},
{-32'd15172, 32'd6814, -32'd2347, 32'd5693},
{-32'd5137, -32'd11829, -32'd6, -32'd6053},
{-32'd16851, -32'd2497, -32'd9039, 32'd4062},
{32'd5360, 32'd14962, -32'd11427, 32'd1848},
{32'd12472, 32'd1846, 32'd3707, -32'd618},
{-32'd5509, -32'd4226, 32'd2103, -32'd2},
{-32'd12117, -32'd4812, 32'd13485, -32'd3628},
{-32'd7709, -32'd5116, -32'd4580, 32'd1172},
{-32'd7773, -32'd7896, 32'd6265, -32'd4381},
{32'd10481, -32'd10851, -32'd3727, 32'd6601},
{32'd2438, 32'd11656, -32'd11158, 32'd11257},
{32'd14083, -32'd7080, -32'd4115, -32'd5569},
{-32'd3789, 32'd14307, 32'd9950, -32'd11919},
{-32'd4336, 32'd7181, -32'd427, -32'd3690},
{32'd3699, 32'd6255, -32'd1797, 32'd13991},
{-32'd6069, 32'd10251, 32'd10058, 32'd1250},
{32'd996, 32'd3242, 32'd32, -32'd3244},
{32'd3919, 32'd1019, -32'd2775, -32'd162},
{32'd9599, -32'd7413, 32'd9573, -32'd8757},
{32'd12376, -32'd11497, -32'd6613, 32'd11167},
{-32'd6244, -32'd359, 32'd781, -32'd2507},
{32'd4630, 32'd7811, -32'd4475, -32'd8742},
{-32'd10076, -32'd4722, 32'd11743, -32'd2943},
{-32'd1804, 32'd8469, 32'd5195, -32'd3229},
{32'd88, 32'd11305, -32'd10088, -32'd7148},
{-32'd8421, -32'd8126, -32'd3165, -32'd1076},
{-32'd8081, 32'd4915, -32'd113, 32'd7479},
{32'd23837, 32'd13160, -32'd4913, 32'd752},
{32'd2590, -32'd10227, -32'd14738, 32'd919},
{32'd17195, 32'd6641, 32'd8174, -32'd6464},
{32'd3202, -32'd3176, 32'd5445, -32'd11183},
{-32'd3057, 32'd6161, -32'd1255, 32'd6875},
{32'd5735, -32'd2277, -32'd13472, 32'd5233},
{-32'd7184, 32'd15401, 32'd1722, -32'd3437},
{-32'd1048, 32'd2484, 32'd11829, -32'd14695},
{32'd2232, 32'd19809, -32'd431, 32'd3214},
{-32'd9141, 32'd9589, 32'd5808, 32'd5311},
{32'd6038, -32'd12002, -32'd2756, 32'd7513},
{-32'd2032, -32'd1094, 32'd5255, -32'd5088},
{32'd5590, -32'd1515, 32'd4861, 32'd15025},
{32'd3244, -32'd1479, -32'd5900, -32'd3683},
{-32'd3252, 32'd1420, -32'd7295, 32'd1500},
{-32'd5098, 32'd7013, 32'd5567, -32'd9710},
{-32'd4488, 32'd5671, -32'd7398, -32'd4067},
{32'd4699, 32'd1787, 32'd7886, -32'd7370},
{32'd9517, -32'd5411, -32'd904, -32'd313},
{32'd1783, -32'd11928, -32'd4877, -32'd9735},
{-32'd206, 32'd269, -32'd1939, -32'd20441},
{-32'd10975, -32'd5371, -32'd11428, -32'd3592},
{-32'd1229, 32'd1945, 32'd1418, -32'd254},
{32'd8559, 32'd8139, -32'd2912, 32'd5851},
{-32'd2997, -32'd14579, 32'd1480, -32'd3715},
{-32'd3091, -32'd5232, 32'd4761, -32'd5193},
{32'd456, -32'd5218, 32'd15777, -32'd6726},
{-32'd23302, 32'd6836, -32'd1125, 32'd287},
{-32'd1697, -32'd3094, -32'd4613, 32'd1665},
{32'd11281, -32'd8120, -32'd9113, -32'd7996},
{-32'd6151, -32'd5218, 32'd5875, -32'd4450},
{32'd4880, 32'd8375, -32'd10471, -32'd1009},
{-32'd7428, -32'd14957, 32'd5550, 32'd1132},
{32'd684, 32'd6286, -32'd354, 32'd2547},
{32'd10148, 32'd6681, -32'd2691, 32'd703},
{32'd6468, -32'd10227, 32'd2401, -32'd5312},
{32'd2042, 32'd4729, 32'd5080, -32'd10865},
{-32'd4729, 32'd167, -32'd1286, 32'd14077},
{32'd1413, 32'd5149, 32'd1072, -32'd8875},
{-32'd8081, -32'd2295, -32'd1252, -32'd2297},
{-32'd2646, -32'd11546, 32'd5241, -32'd10025},
{32'd6372, -32'd1445, 32'd2484, -32'd1472},
{32'd2656, 32'd5336, 32'd9366, -32'd2996},
{-32'd80, 32'd9885, 32'd4944, 32'd22449},
{32'd6947, -32'd8060, -32'd348, -32'd3588},
{32'd12441, -32'd14271, -32'd3902, -32'd798},
{-32'd796, 32'd8948, -32'd4120, 32'd3554},
{-32'd2269, -32'd2530, -32'd9734, 32'd12917},
{32'd4589, -32'd4516, -32'd2665, -32'd9024},
{-32'd8015, 32'd8831, -32'd2384, -32'd2560},
{-32'd875, 32'd10889, -32'd7688, 32'd4519},
{-32'd10336, 32'd9615, -32'd1278, 32'd11043},
{32'd7195, 32'd21818, 32'd2735, -32'd4929},
{32'd11665, 32'd698, 32'd7981, -32'd4294},
{32'd14915, 32'd8014, -32'd6041, -32'd1448},
{-32'd6291, 32'd3169, 32'd3860, 32'd7801},
{32'd5226, 32'd5969, -32'd514, -32'd4760},
{32'd637, -32'd99, 32'd9464, -32'd7811},
{32'd19445, 32'd7994, 32'd5113, 32'd3505},
{-32'd7278, -32'd3975, -32'd832, 32'd2183},
{32'd16914, -32'd3561, 32'd5232, 32'd640},
{32'd11702, 32'd1503, -32'd8887, 32'd3853},
{-32'd1061, -32'd2452, -32'd268, -32'd12768},
{32'd1737, -32'd4812, -32'd6572, 32'd1220},
{-32'd10161, 32'd1452, 32'd12316, 32'd453},
{-32'd5937, 32'd13014, 32'd8447, 32'd15471},
{-32'd9514, -32'd13176, -32'd11748, 32'd1485},
{-32'd3694, -32'd3972, 32'd8874, -32'd324},
{-32'd4325, -32'd13075, 32'd9781, -32'd3925},
{-32'd10619, -32'd6099, -32'd1458, -32'd7749},
{-32'd14632, -32'd22057, -32'd951, -32'd10402},
{32'd2413, -32'd10679, 32'd4791, 32'd2193},
{32'd4132, -32'd3191, -32'd14051, 32'd3505},
{-32'd10247, -32'd1936, 32'd10211, 32'd216},
{-32'd111, -32'd1018, -32'd10354, 32'd3188},
{-32'd5828, 32'd12158, 32'd1980, -32'd849},
{-32'd1499, -32'd14710, 32'd8051, -32'd3580},
{32'd10735, 32'd918, 32'd2118, 32'd3167},
{-32'd14204, -32'd4859, -32'd380, 32'd16083},
{-32'd5556, -32'd7161, 32'd8842, -32'd15429},
{-32'd8476, -32'd1202, -32'd19341, 32'd15145},
{-32'd2008, 32'd6519, 32'd1979, 32'd406},
{32'd2344, -32'd6664, 32'd5072, 32'd8360},
{32'd14514, -32'd6899, 32'd225, 32'd2886},
{-32'd5317, -32'd9281, -32'd7365, -32'd7857},
{32'd7315, -32'd3845, -32'd1419, -32'd643},
{-32'd3082, -32'd1234, -32'd2022, 32'd4612},
{32'd12994, -32'd7030, -32'd11116, 32'd11770},
{32'd3865, 32'd22972, -32'd536, 32'd12026},
{-32'd2393, -32'd6177, -32'd3393, -32'd2820},
{32'd4860, -32'd2057, 32'd790, -32'd2597},
{32'd13572, -32'd7709, -32'd2558, -32'd9749},
{-32'd7504, 32'd16052, 32'd1054, -32'd815},
{32'd991, -32'd766, 32'd4354, -32'd7062},
{-32'd4296, 32'd3262, 32'd7187, 32'd4287},
{-32'd7760, 32'd5735, 32'd7867, 32'd2843},
{-32'd5750, 32'd248, 32'd4971, -32'd2779},
{32'd4829, -32'd2863, -32'd184, -32'd6108},
{32'd9151, -32'd5814, 32'd6659, -32'd2121},
{-32'd3386, -32'd9221, -32'd396, 32'd6506},
{32'd15414, 32'd3364, -32'd5603, -32'd685},
{32'd5591, 32'd5015, -32'd12584, -32'd6095},
{-32'd2012, -32'd5197, -32'd11312, 32'd4652},
{-32'd14339, 32'd14814, 32'd2245, 32'd4098},
{32'd2826, 32'd4793, -32'd3822, 32'd12344},
{32'd8937, -32'd10868, -32'd2689, -32'd2355},
{-32'd2518, -32'd14251, 32'd10160, -32'd8},
{32'd2446, 32'd6500, -32'd10316, 32'd1210},
{-32'd5619, 32'd10736, -32'd8557, 32'd17261},
{-32'd6156, 32'd9848, -32'd2079, 32'd3373},
{-32'd4467, 32'd6454, 32'd3783, -32'd3106},
{32'd3138, 32'd5105, 32'd2226, -32'd6422},
{-32'd7924, -32'd4437, -32'd2369, 32'd2880},
{-32'd3499, -32'd3096, -32'd3145, -32'd6335},
{-32'd13408, 32'd20198, -32'd8304, 32'd6232},
{32'd6699, -32'd3872, 32'd2147, 32'd4434},
{32'd11077, -32'd4233, -32'd2978, 32'd691},
{32'd3384, 32'd11785, -32'd3224, 32'd3527},
{-32'd5402, -32'd711, 32'd12498, -32'd13720},
{-32'd5104, 32'd1624, -32'd10046, 32'd6916},
{-32'd13435, -32'd15845, 32'd4510, 32'd1534},
{32'd4129, -32'd10410, 32'd2737, -32'd7191},
{-32'd6375, -32'd9805, 32'd4642, 32'd11922},
{32'd14620, 32'd13305, -32'd6944, -32'd1083},
{-32'd8120, 32'd1879, 32'd12633, 32'd373},
{-32'd180, -32'd14747, -32'd1789, 32'd9286},
{32'd2806, -32'd7350, -32'd2085, 32'd3204},
{32'd934, -32'd5251, -32'd6412, 32'd11937},
{32'd6122, 32'd7540, -32'd2129, -32'd14993},
{32'd9715, -32'd2260, 32'd858, 32'd1727},
{-32'd2226, 32'd4383, -32'd2358, 32'd5651},
{32'd9442, -32'd7935, -32'd6944, 32'd16241},
{-32'd2590, -32'd4736, -32'd11909, 32'd4232},
{32'd5451, -32'd15109, -32'd1842, 32'd2390},
{32'd5695, 32'd4509, 32'd1053, -32'd3512},
{32'd1819, 32'd16235, -32'd6670, -32'd10166},
{-32'd839, 32'd5753, -32'd2293, 32'd5412},
{-32'd8633, 32'd14146, 32'd9363, -32'd5551},
{-32'd3830, -32'd2226, 32'd9285, 32'd14618}
},
{{32'd14824, 32'd9736, 32'd6734, -32'd7276},
{-32'd23752, -32'd5532, 32'd5937, 32'd1916},
{-32'd7965, 32'd4409, 32'd8485, 32'd2244},
{32'd206, 32'd2313, -32'd399, -32'd1759},
{-32'd888, 32'd19305, 32'd17342, 32'd17108},
{-32'd4820, -32'd4014, -32'd11711, 32'd11866},
{32'd9956, -32'd2294, 32'd8935, -32'd11201},
{-32'd4833, 32'd3903, -32'd1026, -32'd3045},
{-32'd18093, 32'd1528, 32'd7436, 32'd3007},
{32'd4105, 32'd9463, -32'd2191, 32'd2259},
{-32'd6154, -32'd1458, -32'd9204, 32'd2318},
{32'd14030, -32'd1855, 32'd3363, -32'd320},
{32'd3588, 32'd1996, -32'd2604, -32'd7707},
{32'd5966, -32'd4257, -32'd6193, -32'd3554},
{-32'd4479, -32'd6064, -32'd3869, -32'd695},
{32'd10039, -32'd8697, 32'd1162, -32'd5239},
{32'd14317, 32'd17534, 32'd13284, 32'd1310},
{-32'd1392, 32'd1260, -32'd11905, -32'd5927},
{-32'd14095, 32'd5810, -32'd12125, -32'd6623},
{32'd5805, 32'd2433, 32'd11131, -32'd983},
{-32'd6839, -32'd5048, 32'd9280, 32'd4008},
{-32'd9031, 32'd5203, -32'd1366, -32'd2666},
{-32'd14743, -32'd3310, 32'd9965, 32'd3961},
{-32'd6741, -32'd1427, 32'd542, 32'd2983},
{32'd743, 32'd15201, 32'd969, 32'd3703},
{32'd6270, 32'd7435, -32'd6430, -32'd7645},
{-32'd3868, -32'd39, -32'd1724, -32'd7718},
{-32'd17333, 32'd8567, 32'd6695, 32'd9585},
{32'd8058, -32'd4766, -32'd2110, -32'd13568},
{-32'd2235, -32'd4252, -32'd5000, -32'd7654},
{-32'd1637, -32'd19940, 32'd5847, 32'd4698},
{-32'd4120, -32'd6350, -32'd3387, -32'd1844},
{32'd14667, 32'd3863, -32'd2406, -32'd2242},
{32'd5352, 32'd2316, 32'd7942, 32'd1549},
{32'd9633, 32'd13934, 32'd2234, -32'd712},
{-32'd5841, -32'd3028, -32'd3300, -32'd17333},
{-32'd6160, 32'd13322, -32'd7836, 32'd17502},
{-32'd4152, -32'd1351, -32'd1377, -32'd1844},
{32'd16171, -32'd9431, 32'd9001, -32'd872},
{32'd4852, 32'd6318, 32'd524, 32'd1957},
{32'd4828, 32'd13624, -32'd3660, -32'd2154},
{32'd3064, 32'd3524, -32'd2026, -32'd9511},
{-32'd40, 32'd12587, 32'd4708, -32'd837},
{32'd1261, 32'd1491, -32'd9649, 32'd1091},
{32'd2705, -32'd4505, -32'd8302, -32'd2582},
{32'd3386, -32'd9432, 32'd4120, 32'd1623},
{-32'd8008, 32'd3046, -32'd4922, -32'd20417},
{32'd5191, 32'd1996, 32'd2922, -32'd2452},
{-32'd3120, 32'd2692, -32'd10264, -32'd11919},
{-32'd4721, -32'd5756, 32'd14323, 32'd7984},
{32'd6611, 32'd2486, -32'd701, 32'd11009},
{32'd3820, 32'd9675, -32'd6404, 32'd101},
{-32'd10455, 32'd5591, 32'd4228, -32'd10416},
{32'd205, 32'd3559, -32'd6636, 32'd3390},
{32'd4407, 32'd5656, 32'd8294, -32'd4261},
{32'd7243, -32'd1733, 32'd83, -32'd1367},
{-32'd4022, 32'd14, -32'd6115, -32'd4221},
{-32'd2259, -32'd11623, 32'd511, -32'd8531},
{32'd1458, 32'd1032, -32'd9605, 32'd886},
{-32'd2821, 32'd9959, 32'd9023, -32'd4250},
{-32'd6376, 32'd14472, 32'd10763, 32'd2227},
{32'd3177, 32'd4011, 32'd9450, -32'd623},
{32'd488, -32'd11529, -32'd7348, -32'd8068},
{32'd3263, 32'd9908, -32'd6375, -32'd2724},
{-32'd1953, 32'd3539, 32'd9087, -32'd1984},
{32'd6129, 32'd10517, 32'd4448, -32'd2765},
{32'd1463, 32'd4859, -32'd2967, 32'd12047},
{-32'd17409, 32'd3181, 32'd3795, 32'd4398},
{32'd3699, -32'd10194, -32'd866, 32'd55},
{32'd6797, 32'd3598, -32'd115, -32'd1863},
{-32'd4567, -32'd12199, 32'd8816, 32'd4396},
{-32'd14327, 32'd16416, -32'd11710, -32'd12352},
{-32'd9334, -32'd4336, 32'd1827, 32'd1159},
{32'd5181, 32'd6717, 32'd7989, 32'd1833},
{32'd14323, 32'd3066, 32'd14401, -32'd8362},
{32'd16596, -32'd686, 32'd2058, 32'd2193},
{32'd12082, -32'd10815, 32'd15497, 32'd2234},
{32'd4097, 32'd2460, -32'd808, -32'd6223},
{32'd6872, -32'd6212, -32'd8046, -32'd910},
{32'd11634, 32'd7111, -32'd4071, 32'd10724},
{32'd4330, 32'd3052, -32'd19108, -32'd8188},
{32'd5491, -32'd1231, 32'd4006, -32'd5283},
{32'd14971, 32'd1084, 32'd5940, 32'd5468},
{32'd20607, -32'd2253, 32'd7506, 32'd7437},
{32'd8956, -32'd1965, -32'd1881, 32'd126},
{-32'd4998, -32'd4464, 32'd3788, -32'd5591},
{32'd7694, 32'd5317, -32'd3917, -32'd3444},
{32'd25, -32'd1845, -32'd1901, -32'd2034},
{32'd11586, -32'd13133, -32'd5411, 32'd6853},
{-32'd8053, -32'd1715, -32'd4461, 32'd3574},
{-32'd2631, 32'd3657, -32'd3087, -32'd7754},
{-32'd29197, -32'd2584, 32'd1436, -32'd2380},
{-32'd9067, 32'd6979, -32'd11275, -32'd5152},
{32'd13500, -32'd1079, 32'd11288, 32'd9942},
{-32'd490, -32'd5872, -32'd5188, -32'd10954},
{-32'd8693, -32'd4506, -32'd10685, 32'd15632},
{32'd4094, 32'd15327, -32'd601, 32'd2812},
{32'd7484, 32'd7264, -32'd11900, -32'd4648},
{32'd3701, 32'd2829, 32'd7748, -32'd3940},
{32'd4179, 32'd12138, -32'd220, -32'd9575},
{-32'd2137, -32'd14001, -32'd9037, -32'd554},
{-32'd1520, -32'd8128, -32'd1082, 32'd3439},
{32'd9618, 32'd6625, -32'd10321, 32'd15859},
{32'd10036, -32'd2767, -32'd1113, 32'd2856},
{32'd9443, 32'd8447, 32'd5094, 32'd4260},
{-32'd8535, -32'd3321, 32'd8547, -32'd2405},
{-32'd586, -32'd1611, -32'd9369, -32'd101},
{32'd5077, 32'd5830, 32'd10993, -32'd145},
{32'd6195, -32'd5174, -32'd4276, 32'd10710},
{-32'd10438, -32'd5972, -32'd5314, 32'd11470},
{-32'd6432, 32'd15961, 32'd1161, 32'd9445},
{32'd21793, 32'd5744, -32'd940, 32'd2262},
{32'd271, 32'd1077, 32'd12365, -32'd2486},
{-32'd5018, 32'd2553, 32'd3985, -32'd3165},
{32'd2632, -32'd6236, 32'd3180, 32'd6015},
{-32'd6818, -32'd82, -32'd2018, 32'd4373},
{32'd4397, 32'd11756, 32'd7048, 32'd2846},
{-32'd21064, 32'd6431, -32'd4100, 32'd7232},
{32'd12759, 32'd20512, -32'd13691, -32'd12287},
{-32'd6273, 32'd19216, 32'd985, -32'd8524},
{-32'd11120, -32'd2206, -32'd3930, -32'd505},
{-32'd5947, 32'd12499, -32'd6711, 32'd4925},
{-32'd2181, 32'd3339, 32'd2717, -32'd3024},
{-32'd12974, -32'd9501, 32'd204, 32'd7801},
{-32'd8872, -32'd4749, 32'd4606, -32'd4589},
{-32'd9670, -32'd4449, 32'd3611, 32'd5096},
{-32'd16738, -32'd3006, -32'd10086, -32'd4975},
{-32'd13293, -32'd8502, 32'd3594, 32'd3783},
{-32'd14550, -32'd5410, -32'd9278, 32'd2071},
{32'd14164, -32'd8827, 32'd25603, 32'd3015},
{-32'd3979, 32'd12041, 32'd3890, -32'd2728},
{32'd7473, -32'd4714, -32'd3140, -32'd8854},
{32'd10236, -32'd15263, 32'd3031, 32'd9828},
{-32'd2623, 32'd8234, -32'd16782, -32'd9069},
{-32'd11422, -32'd8712, -32'd2836, 32'd2188},
{32'd3024, -32'd6399, 32'd4369, -32'd2703},
{32'd3149, 32'd5229, 32'd6506, 32'd9923},
{-32'd9445, -32'd12559, 32'd5218, 32'd9776},
{32'd3785, 32'd3486, 32'd4580, -32'd15198},
{32'd3357, -32'd9681, 32'd4443, -32'd11499},
{-32'd39, 32'd10762, 32'd881, 32'd1509},
{32'd9941, -32'd4266, -32'd11189, 32'd3274},
{-32'd5799, 32'd14469, 32'd6835, -32'd7069},
{-32'd8820, -32'd6031, 32'd18602, -32'd5750},
{32'd156, 32'd16935, 32'd5250, 32'd14766},
{-32'd7355, 32'd5992, 32'd1171, 32'd9996},
{32'd1391, -32'd6583, 32'd3508, 32'd6815},
{32'd4524, 32'd2030, 32'd6043, -32'd3036},
{32'd2928, -32'd5755, -32'd7185, -32'd3457},
{-32'd3306, -32'd8998, -32'd6607, 32'd5644},
{-32'd1366, -32'd3547, 32'd801, 32'd4152},
{32'd9625, 32'd12557, 32'd10118, 32'd1699},
{-32'd2693, -32'd6426, -32'd7471, 32'd2101},
{32'd16396, 32'd6390, 32'd5819, -32'd667},
{-32'd5647, 32'd772, -32'd8138, -32'd2647},
{32'd4794, -32'd7197, -32'd9087, 32'd663},
{32'd12014, -32'd11982, -32'd8077, -32'd13077},
{32'd10101, 32'd827, -32'd5021, 32'd1904},
{32'd4155, 32'd10937, 32'd4973, -32'd6369},
{32'd10052, -32'd10907, -32'd5471, -32'd10617},
{-32'd6406, -32'd11963, -32'd9634, 32'd10487},
{-32'd2076, 32'd6988, -32'd2576, -32'd272},
{-32'd5227, 32'd558, 32'd11146, -32'd3886},
{32'd2574, 32'd6589, 32'd19406, 32'd4105},
{-32'd3857, 32'd1305, 32'd631, -32'd8224},
{-32'd4045, -32'd8590, -32'd1278, 32'd12911},
{32'd2779, -32'd1907, -32'd13945, 32'd11751},
{32'd2847, -32'd9947, 32'd3868, 32'd4720},
{32'd4812, -32'd474, 32'd10606, -32'd374},
{32'd6606, 32'd329, 32'd2330, -32'd6104},
{32'd1251, -32'd2854, -32'd21844, 32'd1502},
{-32'd4119, -32'd2126, -32'd12411, 32'd892},
{32'd4303, 32'd8120, -32'd5224, 32'd763},
{-32'd7278, 32'd6197, -32'd6477, 32'd12530},
{32'd8827, -32'd939, 32'd9092, -32'd5643},
{32'd6627, 32'd6548, -32'd4575, -32'd622},
{32'd3034, 32'd1467, -32'd3763, 32'd13044},
{-32'd4460, -32'd8883, 32'd1227, -32'd1675},
{-32'd3865, 32'd5612, -32'd1366, -32'd3278},
{-32'd2597, 32'd965, -32'd5205, 32'd4213},
{32'd7988, 32'd3160, 32'd7986, 32'd4032},
{32'd3288, -32'd5771, 32'd2493, 32'd4057},
{-32'd9550, -32'd8107, 32'd2947, -32'd2778},
{-32'd10081, 32'd1169, 32'd4325, -32'd931},
{32'd1478, 32'd6029, -32'd10050, 32'd9214},
{32'd3887, -32'd532, 32'd6793, -32'd4279},
{32'd3191, 32'd6335, 32'd5326, -32'd17415},
{-32'd3064, -32'd647, 32'd5249, -32'd6924},
{-32'd107, 32'd3138, -32'd17007, 32'd6178},
{32'd5125, 32'd1894, -32'd3423, 32'd1944},
{32'd966, -32'd2217, -32'd11510, -32'd9060},
{-32'd11706, -32'd10920, 32'd1355, -32'd1326},
{-32'd11343, 32'd1116, -32'd12203, 32'd2984},
{-32'd13179, 32'd6388, -32'd11528, 32'd11379},
{-32'd5168, -32'd13553, -32'd1074, 32'd3171},
{-32'd9712, -32'd940, 32'd12558, 32'd1275},
{-32'd13383, -32'd14256, 32'd4276, 32'd5287},
{32'd1511, -32'd1059, 32'd7088, 32'd9934},
{32'd2986, -32'd17923, -32'd8421, 32'd1605},
{-32'd11658, 32'd2365, 32'd4990, 32'd10706},
{-32'd9996, -32'd13355, -32'd3720, 32'd2996},
{-32'd5331, 32'd11377, -32'd3326, 32'd3876},
{32'd4970, 32'd1495, 32'd12046, 32'd3500},
{32'd6561, 32'd2999, -32'd3220, 32'd19689},
{32'd741, 32'd6340, -32'd2252, 32'd509},
{32'd6953, -32'd4813, -32'd887, 32'd500},
{32'd9096, 32'd7125, 32'd12279, 32'd980},
{-32'd5827, 32'd406, 32'd973, 32'd1098},
{32'd10554, 32'd3658, -32'd3959, 32'd445},
{32'd5653, 32'd9926, 32'd2002, -32'd1463},
{-32'd1144, 32'd3139, 32'd4122, -32'd1136},
{32'd1271, -32'd2260, 32'd7981, 32'd4366},
{-32'd11608, -32'd2763, 32'd4104, 32'd5404},
{32'd7845, 32'd1411, -32'd75, 32'd4951},
{-32'd14978, 32'd696, 32'd12277, -32'd880},
{-32'd6252, 32'd4056, 32'd1223, 32'd7715},
{-32'd5340, 32'd3672, -32'd10502, 32'd16247},
{-32'd1462, -32'd6032, 32'd2276, 32'd3885},
{32'd25209, 32'd5212, 32'd10425, 32'd7715},
{32'd2679, -32'd373, -32'd1012, -32'd2861},
{32'd11259, -32'd6190, 32'd1754, 32'd2027},
{-32'd10671, 32'd9729, -32'd4923, -32'd3099},
{-32'd3260, -32'd3997, -32'd3267, -32'd4248},
{32'd12482, 32'd625, -32'd3161, -32'd6395},
{-32'd543, -32'd5723, -32'd8522, -32'd3304},
{32'd9851, -32'd10735, -32'd2548, 32'd14098},
{32'd70, -32'd9907, -32'd9009, 32'd3670},
{-32'd16118, -32'd8677, 32'd7955, -32'd8161},
{-32'd1155, -32'd15254, 32'd1047, 32'd6295},
{-32'd5362, 32'd22963, -32'd10497, -32'd3229},
{-32'd4196, -32'd6846, 32'd98, -32'd1911},
{-32'd4824, -32'd58, -32'd3801, 32'd7620},
{-32'd8569, -32'd6958, -32'd10725, -32'd8266},
{-32'd2402, 32'd11399, 32'd6954, -32'd10113},
{-32'd2177, 32'd2915, -32'd15463, -32'd1694},
{-32'd10134, 32'd2068, -32'd10723, -32'd1863},
{-32'd2639, 32'd1704, -32'd3934, 32'd1323},
{-32'd14233, -32'd3640, -32'd10152, 32'd872},
{32'd15519, -32'd6960, 32'd3572, -32'd3340},
{32'd2545, 32'd4242, 32'd2063, -32'd12544},
{-32'd5301, -32'd4153, -32'd252, -32'd16792},
{32'd5392, 32'd5495, 32'd15787, -32'd14874},
{-32'd13488, -32'd9166, -32'd2519, 32'd6905},
{32'd6284, -32'd6006, -32'd323, 32'd8488},
{32'd10463, 32'd10958, -32'd2884, -32'd640},
{32'd16038, 32'd8616, -32'd3410, 32'd8940},
{32'd8645, -32'd7724, -32'd1885, 32'd1238},
{-32'd5440, -32'd2091, 32'd3230, 32'd3889},
{32'd8734, 32'd6181, -32'd1756, 32'd77},
{32'd15946, 32'd7536, -32'd11321, -32'd1731},
{-32'd2077, -32'd7889, 32'd4006, -32'd12075},
{-32'd13451, 32'd4961, -32'd10279, -32'd4792},
{-32'd2279, -32'd1651, -32'd5489, 32'd3676},
{-32'd2200, -32'd9306, -32'd1776, 32'd8479},
{32'd7980, -32'd3321, 32'd5970, 32'd306},
{32'd2211, 32'd1147, -32'd4497, 32'd11691},
{-32'd3171, 32'd8378, 32'd2174, 32'd9676},
{32'd4763, 32'd16778, 32'd3532, 32'd1721},
{32'd8579, -32'd4812, -32'd11337, 32'd3163},
{32'd343, 32'd11673, 32'd3361, 32'd16640},
{-32'd5630, 32'd1033, -32'd13499, 32'd4677},
{32'd9715, -32'd391, -32'd2589, -32'd7154},
{-32'd8713, -32'd23105, 32'd12729, 32'd676},
{-32'd20454, 32'd732, -32'd2725, 32'd7814},
{-32'd2762, 32'd178, 32'd643, 32'd5357},
{-32'd3845, 32'd1261, 32'd5809, -32'd7425},
{32'd8738, -32'd9131, -32'd7749, -32'd10835},
{-32'd792, -32'd8107, 32'd4098, -32'd2953},
{-32'd1852, -32'd4175, -32'd1845, -32'd10073},
{-32'd3622, 32'd1926, 32'd9894, -32'd6300},
{-32'd8158, 32'd4837, 32'd11077, 32'd4120},
{-32'd15866, 32'd16936, 32'd2893, 32'd5690},
{32'd1735, 32'd7494, 32'd5572, 32'd5602},
{32'd1893, -32'd1728, -32'd6079, -32'd2817},
{32'd10766, 32'd2693, 32'd2764, -32'd1066},
{-32'd5070, -32'd2984, 32'd1611, -32'd2654},
{32'd2203, 32'd16741, 32'd2835, -32'd1480},
{32'd1841, -32'd5709, -32'd12352, -32'd9772},
{-32'd1977, -32'd9563, 32'd2178, 32'd1181},
{-32'd5958, -32'd10379, -32'd7360, 32'd5503},
{32'd1423, 32'd7514, -32'd11564, 32'd4278},
{32'd7599, 32'd5447, 32'd10617, -32'd9507},
{32'd14413, -32'd5728, 32'd10923, -32'd7571},
{-32'd7169, 32'd10674, -32'd3919, 32'd273},
{32'd7638, 32'd1595, 32'd11171, -32'd2183},
{32'd1468, -32'd14117, -32'd5173, 32'd4950},
{-32'd13086, -32'd842, 32'd5782, 32'd6262},
{-32'd2626, 32'd1467, -32'd10977, 32'd2793},
{-32'd4045, 32'd7177, -32'd12054, 32'd1703},
{-32'd4996, -32'd7145, -32'd5573, -32'd400},
{32'd11785, -32'd4483, -32'd11813, -32'd3681},
{-32'd2107, 32'd9691, 32'd11819, -32'd873},
{32'd12091, -32'd8285, -32'd7646, -32'd6069},
{32'd4334, -32'd15649, 32'd9469, -32'd542},
{32'd1314, -32'd526, 32'd7095, 32'd6241},
{32'd9605, 32'd1317, -32'd4079, 32'd3677},
{32'd9775, -32'd8672, 32'd12360, -32'd7199},
{-32'd3558, 32'd5009, -32'd7022, 32'd2812},
{-32'd11847, 32'd10802, -32'd4164, 32'd5878},
{-32'd12948, 32'd9273, -32'd3705, -32'd8544}
},
{{32'd4007, 32'd3040, 32'd7293, -32'd2639},
{32'd2579, 32'd3972, -32'd3561, -32'd2135},
{32'd3386, 32'd5715, 32'd6225, 32'd6720},
{-32'd3712, 32'd654, 32'd9401, -32'd880},
{-32'd2725, 32'd6238, 32'd2793, 32'd9067},
{-32'd4753, -32'd13846, -32'd5377, -32'd7047},
{32'd9822, 32'd3181, 32'd7198, 32'd1952},
{-32'd6533, -32'd4072, 32'd1157, -32'd783},
{32'd14513, -32'd3667, 32'd1974, 32'd4340},
{32'd1955, 32'd11559, 32'd697, 32'd1865},
{32'd6076, 32'd1048, -32'd4330, -32'd5390},
{32'd8251, 32'd7810, 32'd7019, -32'd827},
{32'd219, -32'd3200, -32'd885, -32'd4538},
{-32'd4979, -32'd186, -32'd4272, -32'd4508},
{-32'd762, -32'd10485, 32'd3647, 32'd1807},
{-32'd50, -32'd4441, -32'd7009, 32'd6862},
{-32'd4727, 32'd1971, 32'd7045, -32'd451},
{-32'd6618, -32'd11592, -32'd6260, 32'd3116},
{32'd3633, -32'd1003, 32'd5000, -32'd4765},
{32'd10004, 32'd1109, 32'd8137, 32'd9406},
{32'd6696, 32'd2128, 32'd726, -32'd11692},
{-32'd6964, 32'd333, 32'd1755, 32'd1535},
{-32'd6806, -32'd4227, -32'd1011, -32'd611},
{-32'd9748, -32'd5755, -32'd285, -32'd6996},
{-32'd196, 32'd12036, -32'd5712, -32'd10690},
{32'd3278, -32'd2487, 32'd4339, -32'd8712},
{-32'd1443, -32'd4744, -32'd2706, 32'd610},
{32'd12607, -32'd4268, -32'd5169, -32'd5049},
{-32'd3280, 32'd14712, 32'd5529, -32'd2457},
{-32'd2705, -32'd6443, -32'd428, 32'd659},
{-32'd8312, -32'd7441, 32'd13121, -32'd3739},
{-32'd5418, -32'd7028, -32'd7959, 32'd6826},
{-32'd984, 32'd7376, -32'd4524, 32'd3637},
{-32'd876, -32'd4902, -32'd3360, 32'd951},
{32'd9017, 32'd3521, 32'd3014, 32'd8585},
{32'd4244, -32'd6621, -32'd2855, -32'd10265},
{32'd377, -32'd4327, -32'd7203, 32'd5560},
{-32'd989, 32'd2506, 32'd5284, 32'd2816},
{32'd4327, 32'd9582, -32'd3275, 32'd7518},
{-32'd10705, -32'd9203, -32'd4727, 32'd3232},
{32'd2566, 32'd5852, 32'd2752, -32'd2589},
{-32'd3343, 32'd2766, -32'd4009, 32'd4733},
{32'd4514, -32'd480, -32'd3317, 32'd9970},
{-32'd16364, -32'd1197, -32'd2317, -32'd2166},
{-32'd2564, 32'd7601, -32'd72, -32'd305},
{32'd7716, -32'd5835, 32'd2002, -32'd469},
{-32'd2703, -32'd8507, -32'd7890, -32'd1848},
{-32'd3298, -32'd13880, -32'd699, -32'd1235},
{32'd8317, 32'd2476, 32'd2899, 32'd5218},
{-32'd1077, -32'd2603, 32'd6786, -32'd2221},
{32'd13572, -32'd831, 32'd1770, -32'd1518},
{32'd3504, -32'd933, -32'd1294, -32'd8511},
{32'd563, -32'd307, -32'd1875, -32'd4194},
{-32'd16334, 32'd560, -32'd862, 32'd5229},
{-32'd3979, 32'd8545, -32'd1597, -32'd4351},
{32'd8542, -32'd3269, 32'd386, -32'd11017},
{32'd4223, 32'd2817, 32'd5072, 32'd6428},
{-32'd142, -32'd12233, -32'd1866, 32'd2292},
{32'd837, -32'd12507, -32'd2823, -32'd5795},
{32'd9941, -32'd5539, 32'd1927, -32'd5848},
{32'd12047, 32'd2904, 32'd5329, -32'd5785},
{32'd2955, 32'd5405, -32'd5549, 32'd11265},
{-32'd262, -32'd7407, -32'd4048, 32'd3953},
{-32'd338, 32'd4986, 32'd121, 32'd7438},
{-32'd71, -32'd4752, -32'd2626, -32'd1266},
{32'd6444, 32'd5233, 32'd3805, -32'd4003},
{-32'd1812, -32'd3278, -32'd8555, -32'd1705},
{-32'd3111, -32'd184, -32'd189, 32'd5475},
{-32'd3634, -32'd8507, -32'd6711, -32'd6676},
{32'd6796, -32'd4852, 32'd536, -32'd2235},
{-32'd5678, 32'd5545, -32'd6809, 32'd7212},
{-32'd10089, -32'd4769, -32'd1019, -32'd11417},
{-32'd6862, -32'd3260, -32'd5261, -32'd6647},
{-32'd686, -32'd4733, 32'd4634, -32'd2240},
{32'd17819, 32'd7731, 32'd9627, -32'd7799},
{-32'd7808, 32'd8726, -32'd7997, -32'd3048},
{-32'd3842, 32'd1259, -32'd2841, 32'd4200},
{32'd1382, -32'd5630, 32'd273, -32'd7003},
{-32'd4408, 32'd6668, 32'd2216, 32'd4550},
{-32'd9023, -32'd2793, 32'd8411, -32'd1236},
{32'd4286, 32'd4205, -32'd6069, 32'd3552},
{-32'd13198, -32'd3847, 32'd5689, -32'd3331},
{32'd5340, -32'd2735, 32'd5579, 32'd1946},
{-32'd2896, 32'd7643, 32'd371, 32'd1737},
{-32'd7862, -32'd7738, 32'd2312, -32'd7274},
{-32'd2776, -32'd3595, -32'd5599, -32'd5612},
{32'd11180, 32'd1902, -32'd1200, 32'd9097},
{-32'd6436, 32'd6484, -32'd3717, -32'd2337},
{-32'd12627, 32'd1368, -32'd4591, 32'd6890},
{-32'd11353, 32'd9427, 32'd817, -32'd5379},
{32'd4094, 32'd4975, 32'd5323, -32'd658},
{32'd6672, -32'd2192, 32'd83, -32'd2223},
{-32'd8994, 32'd2349, -32'd6456, -32'd490},
{32'd2831, -32'd1869, -32'd262, 32'd11728},
{32'd4876, -32'd4617, -32'd5362, 32'd4783},
{-32'd4342, 32'd2887, -32'd1158, 32'd3568},
{-32'd1689, 32'd8340, 32'd5027, 32'd8516},
{-32'd10466, -32'd7030, 32'd671, -32'd11008},
{32'd5976, -32'd2104, -32'd1634, 32'd5927},
{32'd3070, 32'd5638, 32'd10073, 32'd8337},
{32'd894, -32'd7740, -32'd10648, 32'd1327},
{-32'd4718, 32'd3463, -32'd9411, -32'd3539},
{-32'd3137, 32'd3485, -32'd4603, 32'd736},
{-32'd8079, 32'd10926, 32'd8899, -32'd979},
{32'd5549, -32'd654, -32'd2994, 32'd3430},
{32'd614, -32'd274, -32'd2784, 32'd5862},
{-32'd2174, -32'd3977, -32'd8185, 32'd1461},
{-32'd2342, -32'd1466, 32'd5818, -32'd4503},
{-32'd4396, 32'd2932, -32'd515, -32'd2057},
{-32'd7472, -32'd11890, 32'd1837, 32'd12342},
{32'd11553, -32'd5169, -32'd6574, -32'd7126},
{-32'd6995, 32'd6267, -32'd9768, 32'd1780},
{32'd296, 32'd693, 32'd1109, 32'd5892},
{32'd1069, 32'd4234, -32'd3753, -32'd3728},
{-32'd3819, 32'd2514, 32'd400, -32'd3409},
{-32'd2917, 32'd4604, 32'd1657, -32'd3702},
{32'd4681, 32'd15867, 32'd3248, -32'd3817},
{32'd1195, -32'd5031, -32'd648, -32'd2809},
{32'd3503, 32'd4730, -32'd4260, 32'd2144},
{32'd11837, -32'd648, 32'd3815, -32'd1080},
{32'd5860, -32'd1054, -32'd335, -32'd1975},
{32'd990, 32'd5429, 32'd6171, -32'd2745},
{-32'd3410, 32'd2424, -32'd5301, -32'd2723},
{32'd7770, -32'd2442, 32'd5545, -32'd201},
{32'd4534, -32'd1627, 32'd1048, 32'd1492},
{-32'd434, 32'd4165, 32'd7142, 32'd6599},
{32'd5850, 32'd4164, -32'd4447, -32'd6893},
{32'd3214, -32'd11257, 32'd4957, 32'd687},
{-32'd3263, -32'd6991, -32'd4321, 32'd1340},
{32'd9894, -32'd1795, 32'd2730, -32'd849},
{-32'd760, 32'd1696, 32'd7791, 32'd2917},
{-32'd7152, 32'd1081, -32'd8702, -32'd4643},
{-32'd4180, -32'd4927, -32'd5105, 32'd4812},
{32'd7968, 32'd6148, -32'd4278, -32'd1936},
{-32'd3464, 32'd3118, 32'd2223, 32'd6665},
{-32'd6412, 32'd2083, -32'd290, -32'd806},
{-32'd8208, 32'd1148, 32'd442, -32'd5548},
{-32'd10458, -32'd2729, 32'd8063, 32'd3509},
{32'd10733, 32'd1753, -32'd5176, 32'd6557},
{32'd5473, 32'd416, -32'd5891, -32'd6816},
{32'd6928, 32'd1297, 32'd6568, -32'd1761},
{-32'd5926, -32'd4971, 32'd950, -32'd5635},
{-32'd4057, 32'd6408, -32'd1377, 32'd520},
{32'd2973, 32'd7530, -32'd2006, -32'd1336},
{32'd6724, 32'd9695, -32'd888, -32'd551},
{32'd3346, 32'd6674, -32'd3271, -32'd1527},
{-32'd973, -32'd8829, 32'd8465, 32'd5445},
{-32'd8682, -32'd2295, -32'd3168, -32'd3167},
{32'd6431, 32'd12020, 32'd10172, 32'd1725},
{-32'd17658, -32'd5989, -32'd3004, -32'd10034},
{-32'd13174, -32'd4387, -32'd5011, -32'd424},
{32'd2587, 32'd16526, 32'd13284, -32'd67},
{32'd5305, -32'd3202, 32'd320, 32'd886},
{-32'd1012, 32'd6254, -32'd4167, 32'd3304},
{-32'd9147, -32'd7042, -32'd4582, -32'd656},
{32'd9399, -32'd6686, 32'd161, 32'd9170},
{-32'd1409, 32'd4205, 32'd7726, -32'd1297},
{-32'd5265, -32'd8887, 32'd4627, -32'd5075},
{-32'd4600, -32'd4179, -32'd1393, 32'd7058},
{-32'd2503, -32'd4580, -32'd2359, 32'd4476},
{-32'd666, -32'd12270, -32'd6004, 32'd4172},
{32'd887, 32'd2448, -32'd168, -32'd5704},
{32'd2710, 32'd4642, -32'd5570, 32'd5213},
{-32'd7939, -32'd4678, 32'd7404, 32'd6776},
{-32'd4343, -32'd5479, 32'd483, 32'd3197},
{32'd7320, -32'd13121, -32'd4026, 32'd2229},
{32'd4982, 32'd781, -32'd4175, 32'd1806},
{-32'd12971, -32'd3632, 32'd305, -32'd6377},
{-32'd9363, -32'd433, 32'd25, -32'd1067},
{32'd1049, -32'd11004, 32'd5888, -32'd1194},
{32'd1373, -32'd3049, -32'd12766, 32'd98},
{32'd11591, -32'd4049, -32'd2230, 32'd6988},
{32'd2175, 32'd797, 32'd7695, 32'd5052},
{32'd2868, 32'd503, -32'd2216, 32'd2819},
{-32'd1215, -32'd4434, -32'd3243, -32'd9022},
{32'd3295, 32'd2783, -32'd8548, -32'd152},
{32'd3428, -32'd2987, -32'd7027, -32'd2434},
{-32'd4157, 32'd256, -32'd1046, -32'd5589},
{-32'd12571, 32'd6106, 32'd8272, 32'd105},
{-32'd7901, -32'd5576, -32'd3870, 32'd406},
{-32'd4802, 32'd2179, 32'd158, -32'd14550},
{-32'd14241, -32'd8666, -32'd6315, 32'd6653},
{32'd735, -32'd5062, 32'd874, -32'd11600},
{-32'd6982, -32'd8619, -32'd4636, 32'd3276},
{-32'd1987, 32'd2287, 32'd1913, 32'd6341},
{32'd3675, -32'd3905, 32'd10345, -32'd2681},
{32'd8733, 32'd2620, 32'd5282, 32'd634},
{-32'd3219, -32'd4147, -32'd541, -32'd3518},
{-32'd1393, -32'd10316, -32'd196, 32'd4891},
{32'd486, 32'd6454, -32'd1310, -32'd5224},
{32'd1535, -32'd2434, -32'd2974, 32'd9628},
{-32'd10962, -32'd6187, -32'd8050, -32'd3154},
{-32'd8820, -32'd14504, -32'd7236, 32'd6485},
{-32'd3262, 32'd10232, -32'd6352, -32'd1922},
{-32'd898, 32'd1329, 32'd2509, -32'd2340},
{-32'd3284, -32'd2295, 32'd6365, -32'd1999},
{-32'd6664, -32'd6401, 32'd1809, 32'd6311},
{-32'd886, -32'd3407, 32'd6857, -32'd12515},
{32'd3352, 32'd869, -32'd426, 32'd6570},
{32'd12045, -32'd9929, 32'd1561, 32'd3240},
{-32'd8094, -32'd10629, -32'd6125, -32'd2218},
{-32'd249, -32'd5053, -32'd8164, -32'd7331},
{32'd4628, 32'd1668, 32'd10642, 32'd4185},
{-32'd2349, -32'd1879, 32'd8437, -32'd3955},
{-32'd3302, 32'd4105, -32'd979, 32'd846},
{32'd950, 32'd7579, -32'd2951, 32'd8368},
{32'd6307, -32'd969, 32'd1405, 32'd3309},
{-32'd3282, -32'd9118, -32'd852, 32'd575},
{-32'd2760, -32'd3051, -32'd3528, -32'd3372},
{-32'd1854, 32'd8164, -32'd7281, 32'd7310},
{32'd8413, -32'd3773, -32'd4411, -32'd9254},
{32'd9234, 32'd6651, 32'd6038, 32'd1877},
{-32'd4108, -32'd7422, 32'd583, -32'd898},
{-32'd6446, -32'd7130, 32'd269, -32'd959},
{-32'd2131, 32'd5847, 32'd942, 32'd1397},
{-32'd13238, 32'd987, -32'd2857, 32'd1410},
{-32'd2027, 32'd1191, -32'd5476, 32'd6087},
{-32'd4269, 32'd1999, 32'd102, -32'd9276},
{-32'd6043, -32'd257, 32'd1168, -32'd3139},
{-32'd319, -32'd2914, 32'd4671, -32'd7471},
{-32'd5524, -32'd3860, 32'd4059, 32'd8732},
{32'd16621, 32'd1094, 32'd810, -32'd5112},
{32'd13450, -32'd3124, 32'd5212, 32'd5977},
{32'd4657, -32'd3695, -32'd9544, -32'd16185},
{32'd3485, -32'd11908, 32'd10344, -32'd5911},
{32'd1733, -32'd275, 32'd1690, 32'd3042},
{-32'd10826, 32'd4015, -32'd6850, 32'd1261},
{32'd542, -32'd10450, -32'd710, -32'd4160},
{32'd9705, 32'd2073, -32'd3346, 32'd2646},
{32'd5642, 32'd3922, 32'd5942, 32'd3480},
{-32'd6129, 32'd2357, -32'd4262, -32'd2869},
{32'd10326, -32'd718, -32'd6817, -32'd3078},
{32'd12298, 32'd1483, 32'd2238, -32'd1665},
{32'd296, -32'd6124, -32'd11702, -32'd5306},
{-32'd3002, -32'd7949, -32'd9938, -32'd11394},
{32'd7514, -32'd4748, -32'd6311, -32'd3128},
{32'd655, -32'd2499, -32'd4054, -32'd1426},
{32'd51, -32'd2253, -32'd429, 32'd4982},
{-32'd2422, -32'd6370, 32'd14565, 32'd6032},
{-32'd1960, 32'd5847, -32'd6378, -32'd5021},
{32'd5928, 32'd4138, 32'd3990, -32'd6100},
{32'd15118, -32'd165, 32'd1102, -32'd5687},
{-32'd420, -32'd5809, -32'd5938, 32'd2369},
{32'd8745, -32'd4919, 32'd4101, 32'd4702},
{32'd5092, 32'd11519, 32'd226, 32'd6341},
{32'd543, 32'd764, 32'd9495, -32'd4331},
{-32'd5794, 32'd1610, 32'd5630, 32'd5581},
{32'd1263, 32'd385, 32'd820, -32'd2000},
{32'd4038, 32'd5742, 32'd1367, -32'd5439},
{32'd3899, 32'd11594, 32'd149, 32'd8725},
{-32'd1985, -32'd7646, -32'd5429, -32'd6494},
{-32'd4352, 32'd2443, -32'd6016, -32'd6633},
{32'd1271, 32'd8702, 32'd972, -32'd4095},
{32'd6873, -32'd7151, -32'd6630, -32'd1459},
{-32'd8687, -32'd2203, -32'd1114, 32'd2259},
{32'd5990, -32'd5639, 32'd708, 32'd5680},
{32'd5985, 32'd1433, -32'd6115, 32'd3147},
{-32'd3396, 32'd4885, 32'd7545, -32'd7290},
{-32'd14937, -32'd5493, -32'd7337, -32'd6368},
{32'd12118, -32'd1322, 32'd3206, 32'd74},
{-32'd11, -32'd1141, -32'd1925, 32'd75},
{-32'd16915, 32'd6854, -32'd2451, 32'd2334},
{-32'd5093, -32'd2735, -32'd683, 32'd8549},
{-32'd3714, -32'd791, -32'd3241, -32'd5388},
{32'd3182, -32'd8100, 32'd1413, -32'd435},
{32'd15536, 32'd709, -32'd2808, 32'd2822},
{-32'd5520, -32'd8286, 32'd8099, -32'd609},
{-32'd576, -32'd4811, 32'd1104, 32'd2167},
{32'd1173, -32'd2569, -32'd6680, -32'd5476},
{-32'd9737, -32'd3978, -32'd5817, 32'd8917},
{32'd1378, -32'd8661, 32'd3863, -32'd2593},
{32'd4609, 32'd1355, 32'd7225, -32'd2369},
{-32'd9359, -32'd433, -32'd10216, 32'd2744},
{32'd1312, 32'd252, -32'd4832, -32'd1397},
{32'd2219, 32'd1302, 32'd704, 32'd356},
{32'd8755, 32'd3044, -32'd706, -32'd1506},
{32'd6674, 32'd8889, 32'd5787, 32'd2386},
{32'd5147, -32'd196, 32'd3044, -32'd1276},
{32'd5714, -32'd2588, -32'd1178, -32'd4671},
{-32'd13624, -32'd366, 32'd3600, 32'd4087},
{32'd5310, -32'd551, 32'd2664, -32'd2408},
{32'd6008, -32'd4186, 32'd4639, 32'd17512},
{32'd6737, 32'd4042, -32'd177, 32'd4503},
{-32'd1753, -32'd4836, 32'd7963, 32'd4401},
{32'd19483, 32'd4370, 32'd2915, -32'd1627},
{-32'd7317, -32'd4822, 32'd138, 32'd283},
{32'd4671, -32'd71, 32'd11394, -32'd952},
{-32'd1502, -32'd9940, -32'd11190, -32'd1841},
{-32'd4230, -32'd3691, -32'd4363, 32'd652},
{-32'd9370, 32'd9935, 32'd3808, 32'd1010},
{-32'd7502, 32'd4215, 32'd8813, 32'd1917},
{-32'd4069, 32'd7702, 32'd11825, -32'd1493},
{32'd7947, 32'd4887, 32'd3666, 32'd7475},
{-32'd13640, 32'd4202, -32'd10332, -32'd7083},
{32'd1216, 32'd4034, -32'd1444, -32'd2776},
{-32'd6126, -32'd7346, -32'd786, 32'd1939},
{32'd3103, 32'd3827, 32'd725, 32'd3519},
{-32'd2068, 32'd7906, 32'd1942, -32'd3298},
{-32'd1549, 32'd10068, 32'd8013, 32'd8075},
{32'd14474, -32'd8278, -32'd327, -32'd1230}
},
{{32'd15900, -32'd4105, -32'd5181, 32'd1602},
{32'd3247, 32'd343, 32'd1627, -32'd3412},
{-32'd5667, 32'd1540, 32'd6908, 32'd2058},
{32'd9466, -32'd4591, 32'd10539, 32'd379},
{32'd8251, 32'd7083, 32'd5560, 32'd4378},
{-32'd9720, -32'd5640, -32'd8906, 32'd1616},
{32'd712, 32'd5433, -32'd1448, 32'd2939},
{-32'd10178, 32'd1569, -32'd5118, -32'd9989},
{32'd2342, 32'd1998, 32'd4342, 32'd4829},
{32'd14300, 32'd5909, 32'd12868, 32'd2377},
{32'd1431, -32'd2671, 32'd528, 32'd8114},
{32'd3719, 32'd6855, 32'd2422, -32'd3336},
{32'd571, 32'd4553, 32'd4487, -32'd4352},
{32'd7905, -32'd9138, 32'd1072, -32'd9820},
{32'd1184, -32'd8421, -32'd4658, -32'd8108},
{-32'd1168, 32'd3454, -32'd1569, -32'd5278},
{-32'd51, 32'd13864, -32'd857, 32'd7759},
{32'd3268, -32'd8684, -32'd10668, 32'd3024},
{32'd4374, 32'd4746, -32'd8290, 32'd2134},
{32'd5814, -32'd2496, -32'd3474, 32'd3478},
{32'd1988, -32'd1628, -32'd1497, 32'd9500},
{-32'd5263, -32'd11204, -32'd5017, 32'd3830},
{32'd6636, 32'd3487, -32'd11114, 32'd1047},
{32'd233, 32'd6372, -32'd8590, -32'd10551},
{-32'd7549, -32'd6680, 32'd7795, 32'd3622},
{-32'd2646, 32'd32, -32'd5060, 32'd4046},
{32'd1346, -32'd2800, -32'd11784, 32'd6724},
{-32'd6670, 32'd4398, 32'd9998, 32'd8245},
{32'd6755, 32'd5326, 32'd3185, 32'd2236},
{32'd2739, -32'd4688, 32'd6801, 32'd4065},
{32'd2644, 32'd3974, -32'd7728, -32'd2257},
{-32'd3425, -32'd5581, -32'd7853, 32'd5499},
{32'd9201, 32'd12065, 32'd10080, 32'd9497},
{-32'd13414, -32'd9208, -32'd2690, -32'd3961},
{32'd6578, 32'd4680, 32'd5118, 32'd2966},
{-32'd2624, -32'd9631, -32'd2681, -32'd10510},
{-32'd1586, 32'd1642, 32'd2640, 32'd1699},
{32'd3368, -32'd13783, 32'd68, -32'd6728},
{32'd2676, 32'd2377, 32'd5450, 32'd5026},
{32'd1639, -32'd3934, 32'd6562, 32'd1183},
{32'd2505, -32'd6266, 32'd10415, -32'd927},
{32'd4789, 32'd84, 32'd2254, 32'd3295},
{32'd1422, 32'd10030, 32'd10695, 32'd551},
{-32'd4768, -32'd3207, 32'd1761, -32'd8883},
{32'd9363, -32'd2947, -32'd1028, -32'd11},
{-32'd6513, -32'd5693, -32'd2854, -32'd42},
{-32'd10213, -32'd7505, -32'd1708, 32'd810},
{-32'd6176, -32'd8741, -32'd10369, -32'd5978},
{-32'd1767, 32'd4347, 32'd2098, -32'd6733},
{32'd6076, -32'd306, -32'd6328, -32'd1418},
{32'd2280, 32'd380, -32'd4921, -32'd1775},
{-32'd574, 32'd942, -32'd6887, -32'd9234},
{32'd3754, 32'd1654, -32'd9885, -32'd349},
{32'd5885, 32'd5671, -32'd2426, 32'd2852},
{32'd5013, -32'd1571, 32'd9743, -32'd2456},
{32'd4123, -32'd10653, -32'd3917, 32'd519},
{32'd5718, -32'd3530, 32'd1825, 32'd5716},
{-32'd2397, -32'd4040, -32'd2096, 32'd867},
{-32'd6664, -32'd1841, -32'd7952, -32'd2730},
{-32'd813, -32'd103, -32'd6555, 32'd4162},
{32'd1818, -32'd6621, -32'd11971, -32'd5912},
{-32'd6918, 32'd796, 32'd9954, 32'd7289},
{-32'd5402, -32'd4333, -32'd4643, -32'd2140},
{-32'd5487, 32'd2008, -32'd4569, -32'd1649},
{-32'd5058, -32'd5068, 32'd8279, -32'd7543},
{32'd9738, -32'd4955, 32'd5299, 32'd5096},
{32'd6416, 32'd8363, -32'd3976, 32'd97},
{32'd2799, 32'd8101, 32'd2173, 32'd1113},
{32'd967, -32'd7818, -32'd9743, -32'd1737},
{32'd3780, -32'd5137, -32'd5026, 32'd935},
{32'd12011, 32'd4530, 32'd5495, 32'd4632},
{-32'd7059, -32'd2124, 32'd9596, 32'd1552},
{-32'd10192, -32'd7285, -32'd12329, 32'd2095},
{-32'd8162, -32'd1639, -32'd1436, 32'd3650},
{32'd7901, -32'd2274, 32'd631, 32'd8809},
{32'd6634, 32'd16912, 32'd1004, -32'd384},
{-32'd629, 32'd14158, 32'd163, -32'd2395},
{-32'd9773, 32'd4329, -32'd12804, 32'd949},
{-32'd1165, 32'd5821, 32'd8162, 32'd935},
{32'd13372, 32'd3123, -32'd1625, 32'd8343},
{32'd4308, 32'd4173, -32'd6267, 32'd599},
{32'd2821, 32'd4522, -32'd3326, 32'd2907},
{-32'd7143, -32'd150, 32'd3432, 32'd2385},
{-32'd2746, -32'd1920, 32'd7478, 32'd2763},
{-32'd1009, 32'd4874, 32'd2359, -32'd10870},
{32'd6560, -32'd607, -32'd3152, 32'd495},
{32'd679, -32'd6900, 32'd13719, 32'd2454},
{-32'd8959, -32'd3930, -32'd6281, -32'd10435},
{-32'd3857, 32'd4335, -32'd1148, 32'd1471},
{32'd2398, -32'd2773, -32'd10407, 32'd1176},
{32'd3395, -32'd5788, 32'd8442, -32'd3304},
{-32'd3074, -32'd1362, -32'd3946, -32'd4756},
{32'd7326, 32'd2516, 32'd5350, 32'd1377},
{32'd11765, 32'd8533, 32'd8319, 32'd1735},
{-32'd829, 32'd11814, 32'd2584, -32'd1695},
{32'd4920, 32'd6282, 32'd4970, -32'd4330},
{32'd5478, 32'd3872, 32'd648, -32'd1171},
{32'd8989, 32'd3736, -32'd727, -32'd3984},
{-32'd5449, 32'd1630, 32'd219, 32'd2492},
{32'd14604, 32'd6148, 32'd10129, -32'd150},
{-32'd831, -32'd4492, 32'd9615, 32'd489},
{-32'd6286, -32'd8677, -32'd11383, -32'd180},
{-32'd3934, 32'd5665, 32'd2260, -32'd1200},
{-32'd344, 32'd2755, -32'd893, -32'd807},
{-32'd5657, 32'd1624, 32'd905, 32'd4897},
{-32'd7364, -32'd5215, -32'd8231, 32'd545},
{-32'd3360, -32'd11376, 32'd54, 32'd5672},
{-32'd1600, -32'd3677, -32'd2205, -32'd7962},
{32'd9841, 32'd5600, 32'd5038, -32'd864},
{-32'd4427, 32'd5093, -32'd11543, 32'd1171},
{-32'd3225, 32'd3752, -32'd176, -32'd3130},
{-32'd4675, 32'd2164, 32'd189, -32'd2058},
{-32'd3426, 32'd4768, 32'd2841, -32'd7591},
{-32'd3958, 32'd1790, 32'd2596, -32'd5784},
{32'd836, 32'd2186, -32'd2181, -32'd2634},
{-32'd1849, -32'd3498, -32'd873, 32'd9000},
{32'd6116, -32'd7617, -32'd7001, 32'd1713},
{32'd8556, -32'd1176, 32'd9458, 32'd1177},
{32'd6383, -32'd2089, 32'd4054, 32'd7463},
{32'd4242, 32'd18551, 32'd7188, 32'd902},
{-32'd391, 32'd4797, 32'd3894, -32'd3854},
{-32'd3537, 32'd12630, 32'd10375, 32'd5328},
{-32'd9476, 32'd2974, -32'd2256, -32'd850},
{-32'd53, -32'd4379, 32'd3696, 32'd5788},
{32'd1596, -32'd525, 32'd2019, -32'd481},
{32'd5956, 32'd10715, 32'd2704, 32'd425},
{-32'd739, 32'd387, -32'd697, 32'd3170},
{-32'd374, -32'd11736, -32'd1647, -32'd3924},
{-32'd14132, 32'd7816, 32'd1733, -32'd7070},
{-32'd6514, 32'd4571, -32'd10127, 32'd6800},
{32'd3524, -32'd7055, -32'd8121, 32'd752},
{-32'd2124, -32'd10853, 32'd1944, -32'd2659},
{-32'd4775, -32'd1295, -32'd7144, -32'd1722},
{-32'd260, -32'd7044, 32'd7550, 32'd2954},
{-32'd7906, 32'd7374, -32'd3236, -32'd2494},
{-32'd7778, 32'd13187, -32'd4797, 32'd4642},
{-32'd4258, 32'd1626, 32'd1605, -32'd946},
{32'd8664, -32'd4725, 32'd3424, -32'd6352},
{-32'd8018, 32'd12277, 32'd3908, 32'd253},
{32'd2192, -32'd5572, -32'd3196, -32'd8404},
{32'd1308, -32'd4315, 32'd502, 32'd8434},
{-32'd11906, -32'd4525, -32'd3513, 32'd3533},
{-32'd7839, -32'd4122, -32'd2297, -32'd254},
{32'd3088, 32'd2340, -32'd2105, -32'd1622},
{32'd8093, 32'd6408, 32'd13819, 32'd3132},
{-32'd1657, 32'd7945, 32'd4062, -32'd5271},
{32'd988, 32'd2993, 32'd2112, -32'd2755},
{-32'd4600, -32'd4341, -32'd231, 32'd1797},
{32'd4813, -32'd2610, -32'd2898, -32'd753},
{-32'd5548, -32'd3200, -32'd2968, 32'd1563},
{-32'd5461, 32'd2747, 32'd798, -32'd698},
{-32'd561, 32'd6083, 32'd7409, 32'd1724},
{-32'd3151, 32'd7652, 32'd2963, -32'd1358},
{32'd6445, -32'd4828, -32'd2073, 32'd793},
{-32'd16528, -32'd6624, -32'd11733, -32'd5887},
{32'd3777, -32'd4718, 32'd5466, 32'd3373},
{32'd1669, -32'd7938, 32'd4776, 32'd7363},
{32'd2531, -32'd842, -32'd19963, 32'd1178},
{-32'd9108, -32'd2720, -32'd9461, -32'd3093},
{32'd5331, 32'd1551, 32'd6583, -32'd8733},
{-32'd5535, -32'd7262, 32'd6313, -32'd4236},
{32'd5275, 32'd7525, 32'd7757, 32'd6423},
{-32'd7646, 32'd4176, -32'd4527, 32'd1878},
{-32'd6434, 32'd7641, 32'd11018, 32'd1319},
{-32'd8474, -32'd2204, -32'd3010, 32'd10552},
{32'd1163, -32'd11161, -32'd3603, -32'd2342},
{32'd11711, -32'd1964, 32'd9896, 32'd1841},
{-32'd10244, -32'd1614, 32'd1163, -32'd5205},
{-32'd3001, -32'd2935, 32'd4262, -32'd10618},
{-32'd8523, -32'd6493, -32'd1287, -32'd926},
{-32'd9859, -32'd4026, -32'd7787, -32'd4505},
{32'd1721, -32'd682, 32'd4061, -32'd4258},
{-32'd2331, -32'd314, 32'd2413, 32'd5299},
{32'd185, 32'd1775, 32'd914, -32'd2693},
{32'd8637, -32'd2229, -32'd15846, 32'd1207},
{32'd5112, 32'd371, 32'd9099, 32'd151},
{32'd6978, 32'd1985, -32'd2577, 32'd10985},
{32'd5222, 32'd5059, -32'd10768, 32'd2070},
{-32'd4358, 32'd3100, -32'd3219, 32'd2694},
{-32'd3223, -32'd363, -32'd225, -32'd4964},
{-32'd10585, 32'd5372, -32'd12145, 32'd5283},
{32'd1899, 32'd1845, -32'd44, 32'd1044},
{-32'd2246, 32'd4939, -32'd1471, -32'd4388},
{-32'd516, 32'd4801, -32'd1657, 32'd1854},
{32'd2001, -32'd87, 32'd5017, 32'd3111},
{32'd2555, 32'd3424, 32'd11464, 32'd5072},
{32'd2680, 32'd5447, 32'd2508, -32'd1395},
{-32'd3284, 32'd1614, 32'd1236, -32'd2131},
{-32'd92, 32'd7049, -32'd2623, 32'd1395},
{-32'd2332, 32'd9137, -32'd517, -32'd7516},
{-32'd1195, -32'd5789, -32'd597, -32'd6291},
{-32'd5737, -32'd7122, -32'd7562, -32'd7694},
{-32'd2326, -32'd5959, -32'd4240, -32'd1542},
{32'd5193, 32'd2861, -32'd4515, 32'd569},
{-32'd5145, -32'd5747, 32'd3209, -32'd5965},
{-32'd917, 32'd5317, -32'd5195, 32'd2149},
{32'd2223, -32'd2621, -32'd6894, 32'd1501},
{32'd2464, 32'd4895, 32'd4437, -32'd475},
{32'd2468, -32'd3056, -32'd2896, 32'd8807},
{32'd4648, 32'd8731, 32'd3724, 32'd1413},
{-32'd6456, -32'd7634, -32'd6851, -32'd4010},
{-32'd1289, 32'd5044, -32'd2297, 32'd8974},
{32'd4444, 32'd8226, 32'd7692, -32'd3427},
{-32'd3950, -32'd6463, 32'd2427, 32'd4901},
{-32'd13433, 32'd5117, 32'd9552, -32'd6046},
{-32'd23, 32'd1665, 32'd7223, 32'd4259},
{32'd499, 32'd1925, 32'd12859, -32'd5286},
{-32'd265, 32'd3885, -32'd3648, -32'd7190},
{32'd3486, 32'd14703, -32'd1792, 32'd3565},
{32'd4598, 32'd7975, 32'd3722, -32'd344},
{32'd7918, 32'd1445, -32'd5391, -32'd7241},
{-32'd467, -32'd8077, 32'd1631, 32'd1038},
{32'd2708, 32'd2272, 32'd657, -32'd2403},
{-32'd2177, 32'd10474, -32'd1867, 32'd965},
{32'd614, 32'd801, -32'd6331, -32'd199},
{32'd5244, 32'd993, -32'd5403, -32'd2665},
{32'd3729, -32'd8353, 32'd5217, -32'd2884},
{-32'd3135, 32'd6285, -32'd4234, 32'd2436},
{-32'd10275, 32'd10285, 32'd4535, -32'd1838},
{32'd7068, 32'd12198, 32'd8804, 32'd2223},
{32'd4899, 32'd5852, 32'd7890, -32'd487},
{32'd1043, -32'd8610, -32'd8154, 32'd1932},
{32'd3324, 32'd13144, -32'd7417, -32'd2334},
{-32'd12289, -32'd3029, -32'd7514, 32'd1860},
{-32'd582, 32'd8417, -32'd12813, -32'd6118},
{32'd1728, 32'd5533, 32'd7347, -32'd939},
{-32'd2203, 32'd1111, 32'd2611, 32'd3214},
{-32'd8556, 32'd2265, -32'd1432, 32'd1044},
{-32'd5093, -32'd1952, 32'd883, -32'd1619},
{-32'd5573, 32'd3481, 32'd4845, 32'd801},
{-32'd727, -32'd3966, -32'd4981, -32'd3139},
{-32'd1238, -32'd6207, -32'd2367, 32'd5838},
{-32'd464, 32'd4613, 32'd498, 32'd3398},
{32'd11272, 32'd11812, 32'd1586, -32'd1101},
{32'd4885, -32'd5143, 32'd9589, -32'd3063},
{32'd742, -32'd3303, 32'd63, -32'd180},
{-32'd5668, -32'd14915, 32'd11197, -32'd2478},
{-32'd4443, -32'd3799, 32'd2911, -32'd2304},
{-32'd1826, -32'd1667, -32'd5811, -32'd346},
{-32'd2407, 32'd5595, -32'd5749, -32'd788},
{-32'd6215, 32'd5831, 32'd11262, 32'd7951},
{32'd3871, 32'd2882, -32'd8273, -32'd6908},
{-32'd3499, 32'd3304, -32'd1380, -32'd1024},
{32'd837, -32'd3768, 32'd4373, -32'd5279},
{32'd6930, 32'd6150, 32'd8894, 32'd5344},
{32'd12132, -32'd11121, -32'd466, 32'd4727},
{-32'd8359, 32'd5580, -32'd1107, -32'd10092},
{32'd7972, -32'd2018, -32'd11331, 32'd1199},
{32'd7800, 32'd4141, 32'd1287, -32'd6379},
{32'd3073, -32'd2841, -32'd635, 32'd7339},
{32'd6266, -32'd5764, -32'd5599, -32'd4832},
{32'd4753, -32'd2496, -32'd6180, 32'd1114},
{-32'd2977, -32'd439, 32'd2731, 32'd3560},
{-32'd3267, -32'd1726, -32'd1736, 32'd6637},
{-32'd6713, -32'd2187, -32'd4882, 32'd280},
{32'd3794, -32'd4894, 32'd3900, 32'd1503},
{32'd5293, 32'd8747, 32'd3228, 32'd2244},
{-32'd4664, -32'd2161, -32'd539, 32'd7996},
{-32'd8785, -32'd15435, 32'd4488, -32'd3481},
{-32'd5841, 32'd11588, 32'd7945, -32'd632},
{32'd6343, -32'd12072, -32'd1629, 32'd2512},
{-32'd4607, 32'd8024, 32'd3672, -32'd5464},
{-32'd866, -32'd3229, -32'd4641, 32'd443},
{-32'd7913, 32'd3777, -32'd7025, -32'd4201},
{32'd3544, 32'd1191, 32'd1949, 32'd11002},
{32'd956, -32'd3543, 32'd3311, 32'd7714},
{32'd826, 32'd894, -32'd1653, 32'd2867},
{32'd9662, 32'd5279, 32'd2331, 32'd270},
{-32'd2520, -32'd1689, 32'd561, -32'd7898},
{-32'd9282, -32'd2082, -32'd5441, -32'd2487},
{-32'd5470, -32'd2809, -32'd8241, 32'd6137},
{-32'd890, -32'd3619, -32'd7921, -32'd1339},
{-32'd4976, -32'd1789, -32'd2961, -32'd1867},
{-32'd3110, -32'd2014, 32'd3704, 32'd2387},
{-32'd2261, -32'd5302, 32'd1778, 32'd13055},
{32'd3822, -32'd1920, -32'd8887, -32'd10145},
{32'd12967, 32'd3670, 32'd12064, 32'd4342},
{-32'd3781, 32'd14120, -32'd4346, -32'd792},
{-32'd5802, 32'd1266, -32'd7894, -32'd1598},
{-32'd9947, 32'd2676, -32'd861, 32'd1228},
{32'd11610, 32'd2358, 32'd4021, 32'd2821},
{32'd7960, 32'd5268, 32'd4088, -32'd5900},
{-32'd342, -32'd39, 32'd3224, 32'd768},
{-32'd356, 32'd412, -32'd6770, 32'd5172},
{32'd6675, 32'd6577, -32'd1617, 32'd7045},
{-32'd13247, -32'd7729, -32'd6067, -32'd5714},
{32'd686, -32'd36, 32'd4772, 32'd7837},
{-32'd2512, 32'd4498, 32'd428, 32'd1776},
{-32'd2724, 32'd2086, 32'd2125, -32'd6868},
{-32'd2167, 32'd3792, 32'd2657, 32'd9384},
{32'd5816, 32'd6947, 32'd4309, -32'd7671},
{32'd8067, 32'd3403, -32'd2044, 32'd2247},
{-32'd4272, -32'd9592, -32'd3752, 32'd1737},
{-32'd6055, 32'd4225, -32'd8890, -32'd4661},
{-32'd9679, -32'd9069, -32'd4021, -32'd5178},
{32'd2786, 32'd2664, 32'd3813, -32'd168},
{-32'd900, -32'd1263, 32'd14189, -32'd2822},
{32'd4584, -32'd7026, 32'd8432, -32'd2372},
{32'd2436, -32'd1666, -32'd70, 32'd2492},
{-32'd900, 32'd1612, -32'd2430, -32'd9055}
},
{{32'd5583, 32'd3623, 32'd7539, -32'd197},
{32'd3486, -32'd8718, -32'd409, 32'd11469},
{-32'd5604, -32'd5138, 32'd4446, -32'd2540},
{32'd13394, 32'd10055, 32'd6219, 32'd3580},
{32'd9514, 32'd5642, -32'd2125, 32'd2174},
{32'd1902, -32'd5910, -32'd3, 32'd10080},
{-32'd165, -32'd14441, 32'd2476, -32'd10451},
{-32'd4089, -32'd7185, 32'd4978, -32'd6985},
{32'd3543, 32'd402, 32'd3690, 32'd3439},
{32'd15993, 32'd6672, 32'd7300, 32'd5989},
{-32'd2287, 32'd9836, 32'd6659, -32'd12320},
{-32'd380, -32'd6359, -32'd1709, 32'd7701},
{-32'd316, -32'd104, 32'd12131, 32'd3102},
{32'd105, 32'd3408, 32'd2564, -32'd8626},
{-32'd949, -32'd2461, 32'd1245, -32'd4727},
{32'd1780, -32'd6515, 32'd1137, 32'd1406},
{-32'd9728, 32'd9261, -32'd425, 32'd642},
{32'd322, 32'd1870, 32'd421, -32'd705},
{-32'd8058, -32'd7021, -32'd7164, -32'd2611},
{-32'd16294, 32'd2794, 32'd382, 32'd3434},
{-32'd5288, -32'd5744, 32'd3177, -32'd11818},
{-32'd1140, -32'd6784, -32'd6089, 32'd5454},
{-32'd3629, -32'd469, -32'd948, -32'd1770},
{-32'd6453, -32'd4612, -32'd1007, -32'd7713},
{32'd8912, 32'd202, 32'd6969, -32'd3112},
{-32'd9453, 32'd924, -32'd5651, 32'd84},
{-32'd6297, -32'd10947, 32'd301, 32'd3541},
{32'd4183, -32'd23, 32'd3306, 32'd6198},
{32'd15696, 32'd15015, 32'd3290, 32'd2520},
{-32'd104, -32'd1573, -32'd4364, -32'd628},
{-32'd1884, 32'd3402, -32'd8068, 32'd15237},
{-32'd5166, -32'd2039, -32'd2167, 32'd2692},
{-32'd2061, 32'd4246, 32'd4566, 32'd2061},
{-32'd3099, -32'd14127, -32'd8897, 32'd393},
{32'd9661, 32'd5033, 32'd5205, 32'd2960},
{-32'd13434, -32'd8873, 32'd2971, -32'd8263},
{32'd8851, 32'd96, -32'd6870, 32'd14291},
{-32'd4147, -32'd3693, -32'd4834, -32'd8555},
{-32'd8081, 32'd7333, -32'd338, 32'd4685},
{-32'd9268, -32'd10720, -32'd4739, -32'd6634},
{-32'd1292, 32'd2907, -32'd10956, 32'd6364},
{-32'd4339, 32'd4061, 32'd4897, -32'd5121},
{32'd5934, 32'd3933, -32'd8964, 32'd2129},
{-32'd2399, -32'd18778, -32'd169, 32'd2315},
{-32'd6296, -32'd13585, -32'd4950, 32'd3170},
{-32'd5608, -32'd5694, -32'd8959, 32'd11669},
{-32'd1658, -32'd14295, -32'd7915, -32'd1512},
{-32'd7932, -32'd7284, -32'd5680, -32'd7889},
{-32'd1089, -32'd6636, 32'd13270, -32'd9242},
{-32'd8413, -32'd9941, -32'd1554, 32'd3464},
{32'd4041, -32'd4362, -32'd436, -32'd6394},
{32'd1377, 32'd2779, 32'd2867, 32'd3479},
{32'd415, 32'd16267, 32'd10133, -32'd4595},
{32'd2128, -32'd3980, -32'd4043, 32'd1616},
{-32'd5130, -32'd47, 32'd13076, 32'd6976},
{-32'd3176, -32'd1555, -32'd5308, 32'd9505},
{-32'd6902, 32'd8064, -32'd603, 32'd1048},
{-32'd618, -32'd5198, -32'd1166, -32'd3816},
{-32'd7587, 32'd3003, -32'd7911, 32'd2183},
{-32'd8706, -32'd7491, -32'd6225, 32'd9914},
{32'd2556, -32'd2848, -32'd2514, 32'd1726},
{-32'd302, 32'd10031, 32'd7542, 32'd3683},
{-32'd2966, -32'd10639, -32'd7224, -32'd27},
{-32'd11246, -32'd801, -32'd3981, 32'd3769},
{32'd991, 32'd6346, 32'd3267, -32'd8752},
{32'd6629, 32'd9823, 32'd9559, -32'd7222},
{-32'd3695, -32'd910, -32'd13415, -32'd3788},
{-32'd3346, -32'd3094, 32'd2191, -32'd4280},
{-32'd17650, -32'd3162, -32'd3365, -32'd5505},
{32'd13369, 32'd2278, 32'd66, -32'd8680},
{-32'd3286, 32'd4354, -32'd7911, 32'd13277},
{-32'd2674, -32'd6193, -32'd1846, 32'd5672},
{-32'd11348, -32'd7719, -32'd7246, -32'd267},
{-32'd9772, 32'd4970, -32'd2911, 32'd2490},
{-32'd8905, 32'd17963, 32'd9847, 32'd4173},
{32'd10061, 32'd6238, -32'd11429, 32'd6069},
{32'd1841, -32'd1580, 32'd3012, -32'd11046},
{-32'd7989, 32'd3111, -32'd10070, -32'd6043},
{32'd15947, -32'd1888, 32'd6291, -32'd11256},
{32'd6114, 32'd4875, 32'd119, 32'd5291},
{32'd7247, 32'd3446, 32'd2118, -32'd3643},
{32'd13720, 32'd9624, 32'd2778, 32'd5573},
{-32'd11305, -32'd3454, -32'd18168, 32'd16078},
{-32'd4342, 32'd7679, -32'd1878, -32'd167},
{32'd11061, -32'd8559, -32'd1580, -32'd10593},
{32'd4507, 32'd1922, -32'd2631, -32'd686},
{-32'd3346, 32'd11857, -32'd872, -32'd3046},
{-32'd14396, -32'd2438, -32'd12579, -32'd37},
{-32'd2166, 32'd8119, 32'd931, -32'd2683},
{-32'd2494, -32'd5015, -32'd2634, 32'd3450},
{32'd5950, -32'd8793, 32'd3472, -32'd6492},
{32'd491, 32'd237, -32'd3095, -32'd19052},
{32'd14150, -32'd5513, 32'd11367, -32'd13910},
{32'd3744, 32'd13129, 32'd8555, 32'd2883},
{32'd3865, 32'd12492, 32'd8649, -32'd798},
{32'd8891, -32'd4524, -32'd5132, -32'd10065},
{32'd56, 32'd6051, -32'd177, -32'd2737},
{32'd10513, -32'd10945, 32'd9993, 32'd5366},
{-32'd4596, 32'd8080, 32'd4633, -32'd4496},
{32'd9174, 32'd2819, 32'd8290, 32'd3828},
{32'd3886, -32'd9077, -32'd9747, 32'd799},
{32'd1578, -32'd5025, 32'd961, 32'd14652},
{32'd6149, -32'd1915, 32'd1029, 32'd6217},
{32'd8824, -32'd8765, -32'd2324, -32'd5425},
{32'd8029, 32'd5714, -32'd8195, -32'd11021},
{-32'd4324, -32'd193, -32'd729, -32'd1226},
{-32'd9257, -32'd2305, 32'd423, 32'd7292},
{32'd2691, -32'd2995, 32'd3107, -32'd493},
{-32'd7930, 32'd3445, 32'd6302, -32'd11133},
{-32'd8219, -32'd5945, -32'd8257, 32'd2009},
{32'd7746, 32'd8709, 32'd1494, -32'd4761},
{32'd3639, -32'd91, -32'd6334, 32'd2208},
{-32'd4268, 32'd4473, -32'd1394, 32'd1367},
{-32'd7535, 32'd4575, 32'd517, 32'd16329},
{-32'd9841, 32'd2848, 32'd163, -32'd5676},
{32'd5038, 32'd3706, -32'd6996, 32'd878},
{32'd3645, -32'd5504, 32'd9558, 32'd4419},
{32'd3940, -32'd8075, 32'd10313, 32'd202},
{32'd7112, -32'd301, 32'd4558, -32'd3314},
{32'd18761, 32'd11775, 32'd17387, 32'd7469},
{32'd1662, -32'd3035, 32'd3532, 32'd4005},
{32'd13520, 32'd22536, 32'd7402, 32'd1599},
{-32'd1664, -32'd4933, 32'd2871, 32'd3349},
{32'd3057, 32'd3706, 32'd2658, -32'd5754},
{-32'd3373, -32'd4411, -32'd4229, -32'd5947},
{-32'd823, 32'd11132, 32'd17171, -32'd2196},
{32'd10413, -32'd8727, 32'd3078, 32'd109},
{-32'd8964, 32'd7858, 32'd6433, -32'd16},
{-32'd277, 32'd4667, -32'd7674, 32'd2502},
{-32'd249, -32'd1163, -32'd7510, 32'd11717},
{32'd4093, -32'd5703, -32'd8737, -32'd2247},
{-32'd12010, -32'd14783, 32'd2539, -32'd8999},
{-32'd4358, -32'd7725, -32'd692, -32'd7707},
{-32'd6259, -32'd1842, 32'd6322, -32'd4355},
{-32'd2246, 32'd9710, -32'd23, 32'd1814},
{32'd3889, 32'd2354, -32'd1386, 32'd14994},
{32'd3747, -32'd10448, -32'd6, 32'd10424},
{-32'd758, -32'd3591, 32'd466, 32'd11015},
{32'd5552, 32'd4112, 32'd6948, -32'd5393},
{-32'd16626, -32'd5140, -32'd9161, 32'd4182},
{-32'd6958, 32'd6664, 32'd8218, -32'd1754},
{32'd2544, 32'd3735, -32'd5715, 32'd7034},
{32'd4128, 32'd4357, 32'd6947, -32'd14920},
{32'd241, -32'd2354, 32'd9802, -32'd2304},
{32'd12916, 32'd6974, 32'd8917, -32'd809},
{-32'd5653, 32'd9449, 32'd1433, -32'd4059},
{-32'd516, 32'd3285, -32'd3649, 32'd1279},
{-32'd8624, -32'd5857, 32'd4016, -32'd1482},
{32'd19909, -32'd131, 32'd4517, 32'd2690},
{-32'd15676, -32'd13145, -32'd9971, 32'd5175},
{-32'd7282, -32'd1870, 32'd927, 32'd126},
{-32'd1936, 32'd130, 32'd1372, 32'd1549},
{32'd9099, -32'd7781, -32'd6591, 32'd5152},
{32'd3358, 32'd592, -32'd8950, 32'd12108},
{-32'd14265, -32'd7903, -32'd16373, -32'd1592},
{32'd2028, 32'd13719, 32'd673, -32'd2115},
{-32'd10474, -32'd10732, -32'd2471, -32'd5412},
{-32'd5923, 32'd1119, 32'd7233, 32'd992},
{-32'd3530, -32'd269, -32'd1850, 32'd627},
{-32'd666, -32'd5977, 32'd6181, 32'd8560},
{-32'd10636, -32'd9808, 32'd6340, -32'd14008},
{32'd10366, 32'd7573, 32'd12618, 32'd9356},
{32'd4758, -32'd2233, -32'd5756, 32'd146},
{32'd2700, 32'd18142, 32'd14669, 32'd382},
{32'd3943, -32'd9153, -32'd2792, 32'd5548},
{-32'd9194, -32'd7874, -32'd3465, -32'd3271},
{-32'd755, 32'd1224, 32'd14162, -32'd5438},
{32'd9568, 32'd9146, 32'd5035, -32'd1908},
{32'd1182, 32'd1314, -32'd5831, 32'd5922},
{-32'd2107, -32'd3596, 32'd1163, -32'd6065},
{32'd506, 32'd759, 32'd6904, -32'd7149},
{-32'd224, -32'd14022, -32'd2942, -32'd5429},
{32'd12374, 32'd2056, 32'd4583, 32'd5236},
{32'd2760, -32'd1912, 32'd3110, -32'd11409},
{32'd9483, -32'd2108, 32'd4016, -32'd9257},
{32'd8927, 32'd4372, -32'd561, 32'd3467},
{32'd9391, -32'd4090, -32'd4909, 32'd672},
{32'd6545, -32'd10493, -32'd5361, 32'd11777},
{32'd4867, 32'd294, 32'd7830, 32'd2838},
{-32'd11309, 32'd1712, -32'd4942, 32'd1430},
{32'd4540, -32'd7698, 32'd5120, 32'd7693},
{32'd703, 32'd1957, -32'd10205, 32'd4741},
{-32'd7929, -32'd1102, -32'd3445, -32'd719},
{-32'd1035, -32'd370, -32'd17050, 32'd13240},
{32'd6122, -32'd7524, 32'd4380, -32'd16422},
{-32'd8497, 32'd5030, -32'd1789, 32'd1247},
{32'd305, -32'd2168, 32'd7291, -32'd4139},
{32'd6232, 32'd4876, 32'd2333, -32'd2309},
{32'd5338, 32'd2052, -32'd1387, -32'd13131},
{-32'd1572, -32'd7719, -32'd4887, 32'd6343},
{-32'd1114, -32'd9508, 32'd482, -32'd11796},
{-32'd6150, -32'd15849, 32'd1657, -32'd9382},
{-32'd2677, -32'd6684, -32'd8802, -32'd10272},
{-32'd4559, 32'd742, -32'd274, -32'd7881},
{32'd6459, 32'd7024, -32'd2519, 32'd6558},
{-32'd1650, -32'd196, -32'd3544, 32'd10660},
{-32'd11019, -32'd10210, -32'd12295, 32'd1018},
{32'd11839, 32'd10592, 32'd794, 32'd10366},
{32'd5485, 32'd2694, -32'd3814, -32'd3661},
{32'd5119, -32'd5000, -32'd1992, 32'd15634},
{-32'd17246, -32'd4350, -32'd7627, -32'd585},
{-32'd1434, 32'd8871, -32'd16328, 32'd1327},
{32'd1484, 32'd8218, -32'd6209, 32'd2479},
{32'd1499, 32'd11891, -32'd1075, -32'd350},
{-32'd3032, 32'd9572, -32'd8302, 32'd1076},
{32'd3311, -32'd939, -32'd16259, -32'd8117},
{32'd5402, 32'd643, 32'd6083, -32'd7997},
{32'd3279, 32'd3288, -32'd5443, -32'd889},
{-32'd5485, -32'd557, -32'd3947, 32'd12288},
{32'd12482, 32'd12731, -32'd587, 32'd10825},
{32'd1811, 32'd4649, 32'd25, 32'd869},
{-32'd2836, -32'd2139, 32'd4146, 32'd4156},
{-32'd8341, -32'd4403, 32'd671, 32'd3887},
{-32'd282, 32'd2581, -32'd1803, 32'd1621},
{-32'd14380, 32'd2714, -32'd10973, -32'd553},
{-32'd1999, -32'd4544, -32'd2513, -32'd9536},
{-32'd7110, -32'd3966, -32'd5766, -32'd6377},
{32'd8784, 32'd1568, 32'd6370, -32'd13040},
{-32'd5858, 32'd10734, 32'd3457, 32'd11817},
{32'd232, 32'd7432, 32'd5517, -32'd2487},
{-32'd6845, -32'd3392, -32'd1087, -32'd105},
{32'd6155, 32'd2115, -32'd8352, -32'd6819},
{32'd4291, 32'd10573, 32'd9880, -32'd4466},
{32'd995, -32'd6225, 32'd1034, 32'd10760},
{-32'd1824, 32'd4611, 32'd2028, 32'd1487},
{-32'd2627, -32'd9537, 32'd3803, -32'd8661},
{-32'd6873, -32'd5513, -32'd3371, -32'd2065},
{-32'd7370, -32'd599, -32'd1426, 32'd2784},
{-32'd226, -32'd7243, -32'd3255, -32'd3445},
{-32'd1171, 32'd8367, 32'd5003, 32'd5807},
{-32'd12942, -32'd18868, -32'd5875, -32'd12074},
{-32'd10938, -32'd7249, -32'd2720, -32'd3883},
{-32'd2553, -32'd419, 32'd7640, 32'd7420},
{32'd2677, 32'd5347, 32'd4627, -32'd1266},
{32'd9737, -32'd8456, -32'd1318, 32'd11352},
{-32'd1716, 32'd8147, -32'd11286, -32'd684},
{32'd4519, -32'd10396, 32'd5156, -32'd4538},
{-32'd73, -32'd3274, -32'd2167, -32'd10632},
{32'd5972, -32'd1086, -32'd4328, 32'd17461},
{32'd6214, -32'd3800, 32'd4136, 32'd15417},
{-32'd11887, 32'd11587, -32'd1918, 32'd7603},
{32'd845, 32'd8897, 32'd5734, 32'd3673},
{32'd2318, -32'd4852, -32'd2287, 32'd13025},
{-32'd6970, 32'd6607, 32'd10567, -32'd7741},
{32'd10408, 32'd12902, 32'd4685, 32'd1198},
{32'd3423, 32'd6578, -32'd3994, -32'd10586},
{32'd6882, -32'd3709, -32'd9854, -32'd3151},
{32'd561, -32'd3059, 32'd925, 32'd8290},
{32'd11795, -32'd920, -32'd17, 32'd7269},
{32'd2266, 32'd11832, -32'd4688, 32'd2991},
{32'd4990, 32'd573, 32'd7029, -32'd14176},
{32'd5900, -32'd914, -32'd205, -32'd906},
{32'd8839, 32'd7222, 32'd1105, 32'd10278},
{-32'd3809, 32'd5435, -32'd1672, -32'd9827},
{-32'd9938, 32'd7913, -32'd4012, -32'd7276},
{32'd851, -32'd781, -32'd5634, 32'd10463},
{32'd3923, 32'd7578, -32'd6751, 32'd1144},
{32'd2984, 32'd8139, 32'd20313, 32'd3567},
{-32'd2254, -32'd13417, -32'd12601, -32'd988},
{-32'd12338, 32'd4196, 32'd82, 32'd7169},
{32'd2370, -32'd5183, 32'd15882, -32'd9746},
{32'd369, 32'd5048, -32'd159, -32'd141},
{32'd8170, 32'd2086, -32'd5038, 32'd236},
{-32'd13112, 32'd10971, -32'd3480, -32'd4993},
{32'd3711, -32'd9432, 32'd246, -32'd6273},
{-32'd2824, 32'd8343, -32'd1578, 32'd18814},
{32'd1359, -32'd4300, 32'd11165, 32'd2343},
{32'd3693, -32'd7207, 32'd11864, 32'd1730},
{-32'd13248, -32'd2580, 32'd4245, -32'd11643},
{-32'd5190, 32'd8451, -32'd7474, -32'd2925},
{-32'd283, 32'd3457, -32'd3106, -32'd5788},
{-32'd2924, 32'd15229, 32'd8387, -32'd8495},
{-32'd2492, -32'd323, -32'd14492, 32'd10443},
{32'd1145, 32'd2602, -32'd7325, 32'd9227},
{-32'd4893, 32'd957, 32'd7360, 32'd8452},
{32'd41, 32'd1764, -32'd2873, 32'd7421},
{32'd13419, 32'd5479, 32'd7093, 32'd3327},
{-32'd2998, 32'd3857, 32'd9503, -32'd6638},
{-32'd5232, -32'd1763, -32'd10173, 32'd7084},
{32'd4483, -32'd12782, 32'd1576, 32'd10014},
{32'd16979, 32'd298, 32'd4880, 32'd3750},
{-32'd7953, 32'd7370, 32'd7263, -32'd6231},
{-32'd2258, 32'd12130, -32'd5159, 32'd4952},
{32'd5113, 32'd12597, 32'd1342, -32'd333},
{-32'd1582, -32'd5946, -32'd753, -32'd175},
{32'd9195, -32'd2498, -32'd6091, -32'd5985},
{-32'd330, 32'd6038, 32'd3546, -32'd5022},
{32'd1781, 32'd6609, -32'd2563, -32'd5900},
{32'd10516, 32'd7189, 32'd2288, -32'd6712},
{32'd11168, 32'd617, 32'd167, -32'd500},
{-32'd1482, 32'd4452, 32'd14025, -32'd2865},
{32'd9494, -32'd3018, 32'd11513, -32'd7714},
{32'd277, -32'd4434, 32'd2353, 32'd8040},
{-32'd5073, -32'd10691, -32'd11016, 32'd2116},
{32'd3816, -32'd6495, -32'd277, 32'd2376},
{-32'd14991, -32'd7993, -32'd710, -32'd4782},
{-32'd4448, 32'd4912, 32'd4150, -32'd12294},
{32'd262, 32'd4270, -32'd1547, 32'd3207},
{-32'd4357, 32'd3302, 32'd5712, -32'd866},
{-32'd5224, -32'd6123, -32'd13961, -32'd1377}
},
{{32'd14675, -32'd8362, 32'd7956, -32'd5566},
{-32'd10427, 32'd4254, -32'd15093, 32'd2272},
{32'd8468, 32'd2497, -32'd12255, 32'd7674},
{32'd2606, -32'd8376, 32'd541, -32'd5451},
{32'd8807, 32'd3835, -32'd1871, 32'd7003},
{32'd3433, -32'd183, -32'd2196, -32'd2050},
{32'd1837, 32'd6354, -32'd811, 32'd7386},
{-32'd5925, -32'd10534, -32'd11559, -32'd5400},
{32'd673, 32'd17710, 32'd14609, 32'd17610},
{32'd507, -32'd3555, 32'd2888, -32'd437},
{-32'd5795, 32'd10375, 32'd1320, -32'd418},
{-32'd5527, -32'd19498, 32'd5720, 32'd10020},
{-32'd2975, -32'd9025, 32'd2059, 32'd5660},
{32'd5970, -32'd18840, -32'd5427, 32'd3122},
{32'd1496, -32'd5571, -32'd9704, -32'd5085},
{-32'd9771, 32'd3319, 32'd771, 32'd4796},
{32'd8957, -32'd2095, 32'd2456, -32'd457},
{-32'd4138, -32'd6169, 32'd2899, -32'd6893},
{32'd9810, 32'd4389, 32'd5234, -32'd9661},
{32'd4191, 32'd1577, 32'd13574, -32'd6811},
{-32'd5753, 32'd7115, 32'd4582, 32'd8195},
{-32'd4079, 32'd11229, 32'd3209, -32'd4503},
{32'd9174, 32'd5542, -32'd2139, -32'd9503},
{-32'd4174, -32'd1336, 32'd3187, -32'd2071},
{32'd7543, -32'd3105, 32'd1182, -32'd764},
{-32'd7719, 32'd3166, -32'd6081, 32'd2278},
{32'd7237, 32'd330, -32'd1063, -32'd5492},
{-32'd2663, -32'd1445, 32'd1973, 32'd1780},
{-32'd3891, -32'd7083, -32'd1265, -32'd5470},
{32'd4118, -32'd916, -32'd10184, 32'd14682},
{32'd622, -32'd14399, -32'd5036, 32'd4166},
{-32'd9034, 32'd476, -32'd3170, -32'd3524},
{32'd1455, -32'd778, -32'd6485, -32'd846},
{-32'd8338, -32'd10834, -32'd3234, -32'd5930},
{32'd1799, -32'd3596, -32'd2032, 32'd2737},
{-32'd7872, 32'd4482, -32'd955, 32'd3890},
{-32'd6793, -32'd11695, -32'd6183, 32'd2342},
{32'd5714, -32'd10899, 32'd14017, -32'd1232},
{-32'd2553, -32'd12687, 32'd7443, -32'd1863},
{32'd79, -32'd4659, -32'd12480, -32'd4586},
{32'd7677, 32'd16486, -32'd3829, -32'd2786},
{-32'd10688, -32'd5673, -32'd3858, -32'd2188},
{32'd4760, 32'd606, 32'd4163, 32'd1793},
{32'd1550, -32'd8189, 32'd767, 32'd6930},
{-32'd3636, -32'd5241, -32'd198, 32'd1490},
{32'd1810, -32'd4844, 32'd7928, 32'd14849},
{-32'd592, 32'd16527, -32'd1461, -32'd12206},
{-32'd5871, -32'd5983, 32'd13355, -32'd457},
{32'd3155, -32'd139, 32'd13394, 32'd10499},
{32'd7089, 32'd920, 32'd6380, -32'd9297},
{32'd8898, 32'd6317, 32'd17268, 32'd8678},
{32'd4796, 32'd1440, 32'd9171, -32'd3762},
{-32'd714, 32'd7117, -32'd3823, 32'd6518},
{-32'd10004, 32'd8957, -32'd13527, -32'd5220},
{32'd14446, -32'd7992, -32'd6705, 32'd2994},
{-32'd10897, 32'd3547, 32'd2303, 32'd3572},
{32'd14464, 32'd13152, 32'd11801, 32'd2634},
{-32'd6155, -32'd3534, -32'd2148, -32'd8272},
{-32'd7440, -32'd3721, -32'd396, 32'd2216},
{32'd558, -32'd9922, -32'd3242, 32'd13596},
{-32'd628, 32'd15935, -32'd2099, 32'd4560},
{-32'd12414, -32'd1790, -32'd5630, -32'd1297},
{-32'd2901, 32'd4835, -32'd12161, -32'd1854},
{-32'd5083, -32'd5974, -32'd214, 32'd5495},
{32'd1635, -32'd6649, 32'd7335, 32'd2553},
{-32'd10157, -32'd3481, 32'd5179, 32'd4892},
{32'd2081, -32'd10310, 32'd7574, -32'd381},
{32'd1496, -32'd5738, 32'd10872, 32'd739},
{32'd118, -32'd7451, 32'd3840, -32'd1120},
{-32'd8197, -32'd5317, -32'd11887, 32'd1894},
{32'd6824, 32'd12521, 32'd10152, 32'd8316},
{-32'd7823, 32'd7928, -32'd8270, 32'd4340},
{-32'd3342, 32'd7601, 32'd3516, 32'd2410},
{-32'd6597, 32'd1548, 32'd11649, 32'd10248},
{32'd553, 32'd7131, 32'd5885, 32'd16227},
{-32'd2484, 32'd911, 32'd701, 32'd4955},
{-32'd1668, -32'd3526, -32'd13155, -32'd15238},
{32'd6699, -32'd267, 32'd1106, -32'd4728},
{-32'd1265, -32'd2871, 32'd8810, 32'd18944},
{-32'd7908, -32'd5040, -32'd7941, -32'd1387},
{32'd7949, -32'd15757, -32'd4281, 32'd6485},
{-32'd907, 32'd14732, 32'd13696, 32'd7844},
{32'd565, 32'd6758, 32'd4886, -32'd5185},
{-32'd2701, 32'd1185, 32'd9545, 32'd6644},
{-32'd1349, 32'd753, -32'd10024, 32'd2202},
{32'd5932, -32'd5078, -32'd3161, 32'd15687},
{32'd2259, -32'd4168, -32'd2716, 32'd1150},
{-32'd7447, -32'd2314, -32'd1620, -32'd10938},
{-32'd10769, 32'd632, 32'd11650, -32'd5455},
{-32'd1605, -32'd7158, -32'd4962, 32'd4223},
{32'd8270, -32'd4810, -32'd1327, -32'd4476},
{-32'd514, 32'd1057, -32'd556, 32'd6058},
{-32'd6127, -32'd6025, 32'd5561, -32'd11510},
{32'd190, 32'd505, 32'd7783, 32'd59},
{-32'd7256, 32'd3609, -32'd3159, -32'd6279},
{-32'd8538, 32'd1904, 32'd2618, -32'd6203},
{32'd18301, -32'd1664, -32'd2700, -32'd4884},
{-32'd3289, 32'd1443, -32'd6644, -32'd12474},
{-32'd21855, 32'd576, 32'd2159, 32'd12350},
{32'd6337, -32'd250, 32'd4979, -32'd11966},
{-32'd4595, 32'd22, 32'd663, -32'd2912},
{32'd3249, -32'd2015, 32'd11318, -32'd1505},
{-32'd5382, 32'd2332, -32'd9275, -32'd10420},
{32'd7869, -32'd11094, 32'd9208, 32'd11287},
{-32'd1154, 32'd14720, 32'd6474, 32'd2257},
{32'd8714, -32'd3359, -32'd11956, -32'd2631},
{-32'd6780, 32'd4808, -32'd2952, 32'd4171},
{32'd5585, -32'd8108, 32'd14636, 32'd10554},
{32'd11581, 32'd1580, 32'd3457, 32'd6472},
{-32'd15751, 32'd9625, -32'd2270, 32'd1451},
{-32'd8673, 32'd17382, 32'd10437, 32'd10953},
{-32'd4090, -32'd5852, -32'd1895, -32'd9754},
{32'd4602, -32'd15387, -32'd3439, 32'd2658},
{32'd1161, 32'd4568, -32'd9409, -32'd1972},
{32'd9809, 32'd8647, -32'd12105, -32'd13174},
{-32'd1404, 32'd4362, 32'd2654, 32'd3198},
{32'd8458, -32'd18327, 32'd11051, -32'd2066},
{32'd2239, 32'd2554, 32'd13732, -32'd13388},
{-32'd10730, 32'd15541, -32'd6399, 32'd1331},
{-32'd6917, 32'd3053, 32'd71, 32'd5943},
{32'd10063, -32'd1372, 32'd9939, -32'd5868},
{-32'd2562, 32'd16162, 32'd1474, 32'd942},
{32'd1479, 32'd1305, 32'd10890, 32'd4252},
{32'd5537, 32'd12415, -32'd2098, -32'd243},
{32'd1161, 32'd4639, -32'd495, 32'd1656},
{32'd6584, -32'd4984, 32'd82, 32'd2692},
{32'd10518, 32'd6284, -32'd423, -32'd5273},
{-32'd10105, 32'd14120, 32'd838, 32'd10490},
{32'd3288, 32'd6298, -32'd3605, -32'd16457},
{-32'd1376, -32'd3492, 32'd3136, 32'd7641},
{32'd6359, 32'd11071, 32'd3826, -32'd7937},
{-32'd5497, -32'd10353, -32'd3800, -32'd11706},
{32'd2723, -32'd17678, -32'd4050, 32'd1892},
{32'd703, 32'd1872, 32'd8010, 32'd12345},
{32'd1546, 32'd12918, 32'd4481, 32'd295},
{-32'd9808, 32'd18399, -32'd6355, 32'd13083},
{-32'd5498, 32'd4197, -32'd12256, -32'd692},
{32'd6287, -32'd6818, -32'd1232, -32'd14782},
{32'd7653, -32'd5530, -32'd6575, -32'd8927},
{32'd17824, -32'd298, -32'd12235, -32'd4567},
{32'd8135, 32'd6881, 32'd6025, 32'd1394},
{32'd2381, -32'd1794, -32'd1757, -32'd6808},
{32'd1976, -32'd11286, 32'd7319, -32'd9849},
{32'd3534, 32'd5179, 32'd5575, 32'd10223},
{32'd6985, -32'd14128, -32'd4908, 32'd6880},
{32'd17571, 32'd12225, 32'd7462, -32'd8566},
{-32'd9383, 32'd3259, 32'd5087, -32'd14261},
{32'd2121, 32'd7517, -32'd3907, 32'd3125},
{32'd7563, -32'd6919, 32'd1696, 32'd3132},
{32'd9908, -32'd2797, -32'd3149, -32'd10102},
{-32'd4800, -32'd10944, -32'd5429, -32'd2798},
{32'd9699, 32'd11309, 32'd18402, -32'd3468},
{32'd5103, 32'd7273, 32'd7650, -32'd2402},
{32'd2676, -32'd7377, -32'd14959, -32'd13513},
{-32'd11785, 32'd8236, -32'd5243, 32'd5545},
{32'd13986, 32'd3861, 32'd4839, -32'd8140},
{32'd519, -32'd13200, -32'd31, 32'd6052},
{32'd6483, -32'd15885, -32'd5798, -32'd1374},
{32'd6291, -32'd3186, 32'd2560, 32'd8395},
{-32'd11273, 32'd9067, -32'd8720, -32'd10248},
{32'd8127, 32'd16980, -32'd944, 32'd7740},
{32'd3892, -32'd8597, -32'd10773, -32'd9097},
{-32'd4399, 32'd14419, -32'd5281, -32'd9827},
{-32'd11946, -32'd2025, -32'd310, 32'd2934},
{-32'd481, -32'd13240, 32'd1373, 32'd4952},
{32'd3089, 32'd8958, 32'd3366, 32'd4215},
{-32'd762, 32'd3646, -32'd232, -32'd7363},
{-32'd19955, -32'd388, -32'd5735, -32'd2295},
{-32'd8275, 32'd11316, -32'd153, 32'd774},
{32'd14990, -32'd10337, 32'd775, 32'd7488},
{-32'd4274, -32'd7058, -32'd9781, -32'd4214},
{-32'd5735, -32'd6028, 32'd4298, 32'd3876},
{-32'd7406, -32'd4725, 32'd2433, 32'd6363},
{-32'd11940, -32'd11619, 32'd5684, -32'd7102},
{-32'd9955, 32'd5804, 32'd5843, 32'd197},
{32'd2789, 32'd4257, -32'd8058, -32'd237},
{32'd977, -32'd13978, 32'd4286, -32'd8250},
{-32'd17635, -32'd1709, 32'd5855, 32'd10995},
{32'd110, -32'd2245, 32'd1859, -32'd370},
{-32'd3136, -32'd2901, 32'd4773, -32'd11941},
{-32'd11584, 32'd1655, 32'd2422, 32'd4006},
{-32'd2282, 32'd3636, 32'd2602, -32'd7408},
{-32'd2108, -32'd712, 32'd2229, -32'd1247},
{32'd12833, -32'd7703, 32'd2750, 32'd2177},
{-32'd1, -32'd9353, -32'd2683, -32'd3830},
{32'd1464, -32'd1651, 32'd3939, 32'd8751},
{32'd5673, -32'd5699, 32'd1560, 32'd4478},
{32'd9739, -32'd587, 32'd3504, -32'd1569},
{-32'd12987, 32'd2812, 32'd4868, 32'd12223},
{32'd110, 32'd5114, -32'd12108, -32'd13212},
{-32'd6081, -32'd7891, -32'd13970, -32'd4222},
{-32'd1235, 32'd7598, -32'd4839, -32'd11938},
{-32'd4005, -32'd2094, -32'd3084, 32'd9572},
{32'd4, -32'd1972, -32'd3677, 32'd1898},
{-32'd12793, -32'd1048, 32'd10144, 32'd8974},
{32'd8189, 32'd4136, 32'd2744, -32'd6959},
{-32'd9618, -32'd6605, 32'd15031, -32'd9535},
{32'd17011, 32'd2950, 32'd2300, 32'd12158},
{-32'd5907, -32'd1918, 32'd7735, -32'd741},
{32'd2564, -32'd6790, -32'd777, -32'd7660},
{-32'd1750, 32'd7760, 32'd3001, -32'd3815},
{-32'd858, 32'd11360, -32'd540, -32'd8839},
{32'd4863, 32'd11146, 32'd5268, -32'd1525},
{32'd10598, 32'd16713, 32'd9103, 32'd829},
{-32'd14605, 32'd1656, -32'd12832, -32'd4480},
{-32'd19495, -32'd3879, 32'd8640, -32'd9360},
{32'd2320, 32'd11017, 32'd12052, -32'd3243},
{32'd2948, -32'd7220, 32'd3015, -32'd1630},
{-32'd15219, 32'd1998, -32'd1678, 32'd2073},
{-32'd7669, 32'd4744, 32'd13903, -32'd12417},
{-32'd11576, 32'd7692, -32'd17388, 32'd11812},
{32'd8546, -32'd15863, 32'd11778, 32'd7452},
{32'd149, 32'd505, -32'd4961, 32'd3752},
{32'd1979, 32'd4372, 32'd5515, -32'd9109},
{32'd11152, 32'd6064, -32'd4914, -32'd12499},
{32'd17347, -32'd8860, 32'd4622, -32'd1828},
{-32'd11747, -32'd3718, -32'd7087, 32'd8838},
{-32'd1530, -32'd1321, 32'd14228, 32'd1380},
{32'd14485, -32'd19154, 32'd16445, -32'd1452},
{-32'd5575, 32'd8862, -32'd11592, 32'd3284},
{-32'd6006, 32'd320, 32'd3269, -32'd7539},
{32'd5036, 32'd11535, 32'd3830, 32'd4786},
{32'd7599, -32'd6007, -32'd3402, 32'd4254},
{32'd6087, -32'd2458, 32'd6059, 32'd483},
{-32'd12554, -32'd2297, -32'd4249, -32'd15137},
{-32'd16626, -32'd7444, -32'd11148, 32'd10834},
{-32'd136, 32'd1919, 32'd8545, 32'd8211},
{-32'd6234, -32'd8140, -32'd2042, -32'd283},
{32'd10196, -32'd2884, 32'd7467, -32'd12523},
{32'd6275, 32'd10834, -32'd8236, -32'd2510},
{-32'd58, 32'd4594, 32'd1790, -32'd2990},
{-32'd5417, 32'd2432, 32'd11547, 32'd8069},
{-32'd10630, 32'd3473, -32'd2693, 32'd2429},
{32'd5608, 32'd15555, -32'd15165, -32'd10472},
{32'd2469, -32'd4308, -32'd14383, -32'd1806},
{-32'd804, 32'd19263, -32'd2624, -32'd2446},
{32'd4466, -32'd9230, 32'd4285, 32'd1541},
{-32'd3589, 32'd151, 32'd4296, 32'd13811},
{-32'd1610, -32'd5068, 32'd9342, -32'd2553},
{-32'd2827, -32'd3378, -32'd12877, 32'd878},
{32'd5425, 32'd9302, 32'd1782, 32'd6859},
{-32'd4946, -32'd11152, -32'd14680, 32'd4061},
{-32'd3214, -32'd4396, -32'd4136, -32'd3018},
{-32'd6295, -32'd8345, 32'd1865, 32'd11286},
{32'd10456, -32'd1254, 32'd1037, 32'd97},
{-32'd2342, -32'd1171, -32'd7347, -32'd10657},
{-32'd8158, 32'd1549, -32'd58, -32'd10227},
{32'd8192, -32'd4644, 32'd8512, 32'd3088},
{-32'd10977, 32'd849, -32'd1931, -32'd12708},
{32'd5452, -32'd7255, -32'd7245, 32'd19241},
{-32'd5968, 32'd6002, -32'd5727, 32'd5057},
{32'd15141, 32'd8117, -32'd14216, -32'd11065},
{32'd12407, 32'd2605, 32'd2289, -32'd7703},
{32'd7740, 32'd14268, 32'd3887, 32'd10802},
{32'd7051, 32'd13929, 32'd8444, 32'd3652},
{32'd1199, 32'd3959, 32'd4766, 32'd2963},
{32'd2949, -32'd6997, 32'd3152, 32'd1610},
{32'd12421, 32'd4782, -32'd2986, -32'd1972},
{32'd773, 32'd2930, -32'd11246, -32'd20578},
{32'd2207, -32'd9169, 32'd3361, 32'd9474},
{32'd4746, 32'd3200, 32'd13579, 32'd1475},
{-32'd1066, -32'd3844, -32'd10678, 32'd1318},
{-32'd4430, -32'd13610, -32'd2618, 32'd11810},
{-32'd10239, 32'd3938, -32'd7233, -32'd604},
{32'd4615, -32'd9405, 32'd9744, 32'd2582},
{-32'd556, 32'd6472, -32'd2251, -32'd4925},
{32'd3940, -32'd11941, -32'd1819, -32'd3765},
{-32'd14369, -32'd3691, -32'd19000, -32'd6602},
{-32'd744, -32'd1490, -32'd12035, 32'd4122},
{-32'd3586, -32'd6762, 32'd1843, -32'd3933},
{-32'd5183, -32'd11775, 32'd9930, 32'd9247},
{-32'd1328, 32'd80, 32'd3240, 32'd14847},
{-32'd11408, 32'd14613, 32'd5061, 32'd1264},
{-32'd761, -32'd1175, 32'd12750, 32'd7991},
{32'd13953, 32'd14618, 32'd4086, -32'd1273},
{-32'd18379, 32'd8730, -32'd1878, 32'd806},
{32'd1753, -32'd1952, 32'd2695, -32'd1539},
{32'd1978, -32'd9385, 32'd4954, 32'd10068},
{32'd1184, 32'd3607, 32'd2315, 32'd1236},
{-32'd6505, -32'd12276, -32'd12340, -32'd6741},
{-32'd2571, 32'd17645, -32'd2691, -32'd248},
{-32'd714, 32'd3864, 32'd15759, 32'd10357},
{-32'd26, 32'd8338, 32'd10958, 32'd3948},
{-32'd12603, 32'd7890, -32'd1005, 32'd8586},
{32'd17404, -32'd5543, 32'd2355, -32'd8441},
{-32'd3600, 32'd2950, -32'd6007, -32'd2231},
{-32'd1205, 32'd11935, 32'd26188, 32'd448},
{-32'd2298, 32'd3933, 32'd1959, -32'd5432},
{-32'd319, -32'd4087, -32'd4051, 32'd4405},
{-32'd3563, 32'd13110, -32'd8694, -32'd6183},
{-32'd7590, -32'd5510, -32'd5282, 32'd15364},
{32'd11073, 32'd4061, 32'd7609, 32'd4007},
{-32'd2577, -32'd342, 32'd6667, -32'd4664},
{32'd7120, -32'd7390, 32'd3326, -32'd4113},
{32'd2767, 32'd6123, -32'd2228, -32'd9265},
{-32'd2908, -32'd1617, -32'd6446, -32'd545},
{32'd7477, -32'd5573, 32'd2706, -32'd5949},
{32'd11382, 32'd359, 32'd5555, 32'd2062},
{32'd6734, -32'd5066, 32'd6941, 32'd4005},
{32'd12030, 32'd11154, 32'd7086, -32'd11660}
},
{{-32'd1257, 32'd1045, 32'd8594, 32'd1307},
{-32'd3378, -32'd2481, -32'd6511, -32'd11855},
{-32'd5455, -32'd2226, 32'd7466, 32'd2453},
{32'd8560, 32'd7712, 32'd36, -32'd461},
{32'd143, -32'd6834, -32'd9222, 32'd11090},
{-32'd5854, -32'd3882, 32'd4993, -32'd6906},
{-32'd6991, 32'd3913, 32'd861, -32'd3207},
{-32'd5924, 32'd3268, 32'd3521, 32'd4010},
{-32'd8986, -32'd4426, -32'd3896, -32'd3394},
{32'd9341, 32'd14179, 32'd9954, 32'd6341},
{-32'd15522, 32'd5053, 32'd10698, -32'd7396},
{32'd9644, -32'd2594, 32'd2982, -32'd7183},
{32'd5722, -32'd5151, 32'd11368, -32'd2899},
{32'd4377, -32'd2491, -32'd3684, -32'd1105},
{-32'd5708, 32'd703, -32'd8242, -32'd1853},
{-32'd490, 32'd3554, 32'd95, -32'd5117},
{32'd2913, 32'd5855, 32'd10109, 32'd10891},
{-32'd9479, -32'd2146, 32'd2984, 32'd2812},
{32'd13461, 32'd473, -32'd228, -32'd2717},
{32'd990, 32'd2528, -32'd979, 32'd124},
{32'd3951, 32'd8767, -32'd3269, -32'd3289},
{-32'd11344, -32'd5330, 32'd2957, -32'd5826},
{32'd8703, 32'd1013, -32'd47, 32'd1314},
{-32'd62, -32'd13315, 32'd4313, -32'd5152},
{32'd7290, 32'd2423, 32'd8588, 32'd3047},
{-32'd7916, -32'd3339, 32'd2177, 32'd4603},
{-32'd4334, 32'd4423, -32'd1239, -32'd2825},
{-32'd1920, 32'd1685, 32'd9483, 32'd4056},
{-32'd8666, 32'd4450, 32'd420, 32'd2196},
{-32'd12229, -32'd2152, -32'd10614, 32'd2260},
{32'd9539, -32'd820, -32'd5449, -32'd9378},
{-32'd11965, -32'd16756, -32'd10340, -32'd170},
{32'd8080, 32'd1701, 32'd15382, 32'd21452},
{32'd3420, -32'd6519, -32'd4613, 32'd2619},
{32'd6551, 32'd3166, 32'd7251, 32'd2145},
{32'd2605, -32'd12182, -32'd379, 32'd4752},
{32'd2806, -32'd2180, -32'd7804, 32'd4810},
{-32'd6626, -32'd11848, -32'd6164, 32'd2371},
{-32'd5548, 32'd5838, 32'd304, -32'd5415},
{-32'd1000, 32'd11458, -32'd1132, -32'd8707},
{32'd3649, 32'd13312, -32'd10238, -32'd3179},
{-32'd2489, -32'd2193, 32'd12023, 32'd3505},
{32'd1336, 32'd10242, 32'd7323, 32'd7737},
{32'd1724, -32'd2777, -32'd3361, 32'd3413},
{-32'd503, -32'd9565, -32'd418, 32'd82},
{-32'd800, -32'd4758, -32'd468, -32'd9762},
{-32'd3667, -32'd11177, 32'd7048, 32'd6082},
{-32'd5763, -32'd4096, -32'd10013, 32'd713},
{32'd3343, 32'd10051, 32'd11806, 32'd9255},
{32'd305, 32'd1403, 32'd9728, 32'd6912},
{-32'd842, -32'd4407, -32'd985, 32'd2386},
{-32'd1246, -32'd10651, -32'd3707, 32'd174},
{32'd4009, -32'd565, 32'd8149, -32'd1875},
{32'd6489, 32'd3754, -32'd16666, 32'd9262},
{32'd10891, 32'd3594, -32'd272, -32'd1715},
{-32'd3660, 32'd780, -32'd8632, 32'd2002},
{32'd1816, 32'd10523, 32'd7486, 32'd6047},
{-32'd5087, -32'd8573, -32'd8252, -32'd1315},
{32'd1405, 32'd7131, -32'd9254, -32'd7130},
{-32'd2471, -32'd1146, -32'd2456, -32'd10325},
{-32'd5272, -32'd12707, -32'd9122, 32'd2859},
{-32'd8721, 32'd7252, -32'd2343, -32'd280},
{32'd3599, -32'd14023, -32'd2337, -32'd8313},
{-32'd4846, -32'd7650, -32'd7875, -32'd6766},
{32'd1936, 32'd13192, 32'd9685, 32'd11557},
{32'd6001, -32'd1593, 32'd16178, 32'd4422},
{-32'd2502, 32'd748, -32'd11242, -32'd14748},
{32'd1512, -32'd3744, 32'd1552, -32'd5104},
{32'd1259, 32'd9118, -32'd3551, 32'd769},
{32'd3837, 32'd1881, -32'd300, -32'd6064},
{-32'd853, -32'd3387, -32'd8122, -32'd3798},
{-32'd4233, -32'd2171, 32'd18011, -32'd330},
{-32'd13648, -32'd520, -32'd7311, 32'd2452},
{32'd1652, 32'd5279, 32'd9782, 32'd11119},
{-32'd12136, 32'd5529, 32'd5774, 32'd1700},
{32'd938, -32'd8806, -32'd2563, -32'd971},
{32'd5229, -32'd7058, -32'd7037, -32'd7855},
{32'd5471, -32'd7176, -32'd2727, -32'd7514},
{32'd5688, -32'd1228, 32'd6264, 32'd8278},
{-32'd5416, 32'd1906, 32'd8336, -32'd1995},
{32'd4947, 32'd7354, -32'd9522, -32'd6218},
{32'd5758, 32'd11508, 32'd11590, 32'd11610},
{32'd5526, 32'd4564, -32'd12824, -32'd3715},
{-32'd1640, -32'd3551, -32'd2311, -32'd3302},
{-32'd5294, -32'd13436, -32'd9490, 32'd2569},
{32'd4725, -32'd1183, -32'd201, -32'd7090},
{-32'd12197, 32'd2844, 32'd14876, 32'd11024},
{32'd3183, -32'd6169, -32'd3457, -32'd4462},
{-32'd1841, 32'd724, -32'd5526, -32'd3319},
{32'd9339, 32'd2771, -32'd5456, -32'd6381},
{32'd1976, 32'd2803, 32'd11733, -32'd1614},
{32'd2289, -32'd7098, 32'd1110, -32'd10866},
{32'd4365, 32'd606, 32'd6801, 32'd5405},
{32'd4974, 32'd1009, 32'd9637, 32'd560},
{-32'd16145, -32'd4508, 32'd16906, 32'd7773},
{-32'd6089, 32'd4998, -32'd8078, -32'd1696},
{32'd11032, 32'd8017, -32'd4268, 32'd6803},
{-32'd2895, -32'd11780, 32'd1215, 32'd5548},
{-32'd5517, -32'd16404, -32'd5026, 32'd543},
{32'd16320, 32'd3499, -32'd2246, 32'd2119},
{-32'd4225, 32'd5330, 32'd3996, -32'd4452},
{-32'd870, -32'd5580, 32'd5979, -32'd3560},
{-32'd11204, 32'd4108, -32'd5442, -32'd6399},
{32'd9867, 32'd5568, -32'd2070, -32'd100},
{-32'd5213, 32'd9942, 32'd5002, 32'd12679},
{-32'd13048, 32'd8869, -32'd8196, -32'd8461},
{-32'd8813, 32'd3002, 32'd25, -32'd1519},
{32'd9146, -32'd11129, -32'd6093, -32'd1764},
{-32'd965, 32'd10237, -32'd5248, 32'd3331},
{32'd2446, -32'd5129, -32'd6147, -32'd624},
{-32'd5017, 32'd6785, -32'd5599, 32'd4501},
{32'd4605, 32'd4768, -32'd1775, -32'd4787},
{32'd10435, 32'd11010, 32'd4764, -32'd2259},
{-32'd1282, 32'd625, 32'd7439, -32'd6406},
{-32'd1414, 32'd2260, -32'd6782, -32'd1643},
{32'd5881, 32'd6557, -32'd15286, 32'd1344},
{-32'd1825, 32'd6608, 32'd521, 32'd102},
{32'd2600, -32'd3191, 32'd8737, -32'd3436},
{-32'd4610, 32'd12362, -32'd2744, 32'd3346},
{32'd8101, 32'd6390, 32'd20548, 32'd8024},
{32'd13526, -32'd321, -32'd2255, 32'd1444},
{32'd5117, 32'd738, -32'd3813, 32'd6216},
{32'd3326, -32'd3428, 32'd4778, 32'd4176},
{-32'd2963, -32'd1041, -32'd9788, 32'd3478},
{-32'd1413, 32'd7693, -32'd4448, 32'd7003},
{32'd9953, 32'd5995, 32'd4771, 32'd1596},
{32'd899, 32'd11199, -32'd4532, -32'd5367},
{-32'd18445, -32'd203, -32'd4838, 32'd10631},
{-32'd6942, 32'd101, -32'd3798, -32'd2346},
{32'd13738, -32'd15349, 32'd370, -32'd4698},
{32'd945, -32'd14647, 32'd1596, 32'd11303},
{-32'd1988, -32'd6519, -32'd1427, 32'd1633},
{-32'd16520, -32'd3091, -32'd7370, -32'd12670},
{32'd5268, -32'd1082, 32'd6862, 32'd48},
{32'd7387, -32'd7429, -32'd4239, 32'd7892},
{32'd6228, 32'd1505, 32'd8714, -32'd331},
{32'd3636, 32'd1246, 32'd2193, -32'd3079},
{32'd7957, -32'd7415, -32'd14887, -32'd8825},
{32'd6544, 32'd8130, -32'd1759, 32'd2099},
{-32'd2332, -32'd12187, -32'd2350, -32'd4813},
{32'd1228, 32'd1817, 32'd2517, 32'd812},
{-32'd601, 32'd2434, -32'd2378, -32'd3401},
{-32'd1838, -32'd6253, 32'd5125, -32'd403},
{-32'd6809, -32'd3156, 32'd112, 32'd4967},
{32'd6738, -32'd2164, 32'd11314, 32'd7449},
{-32'd5990, 32'd3675, 32'd6428, 32'd3647},
{-32'd11310, -32'd812, 32'd8848, -32'd537},
{-32'd1791, 32'd11526, -32'd5892, -32'd6639},
{32'd7712, -32'd6328, -32'd1046, 32'd188},
{-32'd648, -32'd3006, 32'd6585, -32'd8719},
{-32'd64, -32'd4187, -32'd540, -32'd3686},
{32'd3997, 32'd7124, 32'd9150, 32'd6664},
{32'd3662, -32'd9559, 32'd1871, 32'd8185},
{32'd1113, 32'd622, -32'd8263, -32'd13301},
{-32'd2708, -32'd5492, -32'd10846, -32'd1840},
{32'd142, -32'd1658, -32'd13542, 32'd1932},
{32'd7141, 32'd5903, 32'd6015, 32'd2278},
{-32'd7008, 32'd9371, 32'd5140, 32'd35},
{32'd5510, -32'd7033, 32'd4420, -32'd2070},
{-32'd5398, -32'd9036, -32'd791, 32'd2105},
{-32'd12411, -32'd11617, 32'd6619, 32'd7989},
{32'd8299, -32'd7943, 32'd7782, 32'd5836},
{32'd2388, 32'd918, -32'd25067, -32'd1255},
{-32'd9347, 32'd7255, 32'd3571, 32'd3489},
{32'd7782, 32'd1411, -32'd2632, -32'd10329},
{-32'd4171, 32'd4733, 32'd126, 32'd1948},
{-32'd15242, 32'd9327, 32'd2283, 32'd2318},
{-32'd10556, -32'd7869, -32'd4146, 32'd4782},
{-32'd6079, -32'd716, -32'd8045, -32'd8815},
{-32'd10719, -32'd13790, 32'd12609, 32'd5948},
{-32'd12568, 32'd4417, -32'd13862, -32'd2210},
{32'd2342, -32'd5244, 32'd2268, 32'd15005},
{32'd7903, 32'd14244, 32'd5216, 32'd5546},
{32'd7678, -32'd4036, 32'd9880, -32'd854},
{32'd9952, 32'd3373, -32'd9803, 32'd25},
{32'd8262, -32'd8794, 32'd2144, 32'd3456},
{32'd4946, 32'd14239, 32'd6497, 32'd7348},
{-32'd12481, 32'd9, -32'd9734, -32'd2654},
{32'd6483, -32'd4280, 32'd15291, 32'd9777},
{-32'd12200, 32'd7465, -32'd4007, 32'd371},
{-32'd1067, 32'd3554, 32'd2701, 32'd576},
{32'd4103, 32'd3835, -32'd1043, 32'd2355},
{32'd5052, 32'd4132, -32'd2782, -32'd2925},
{-32'd2876, -32'd1248, 32'd6874, -32'd2991},
{-32'd2618, 32'd7293, 32'd14783, 32'd10748},
{32'd1226, 32'd14272, -32'd4833, 32'd369},
{-32'd1435, -32'd6137, 32'd4605, -32'd6967},
{32'd2590, 32'd4993, 32'd9494, 32'd3263},
{-32'd14342, 32'd1267, -32'd540, -32'd3480},
{32'd896, -32'd1782, -32'd13895, -32'd2739},
{-32'd12470, -32'd10183, -32'd12338, 32'd9232},
{32'd7866, -32'd7415, -32'd12025, 32'd3330},
{32'd584, 32'd19271, -32'd11757, -32'd372},
{-32'd3081, -32'd2643, 32'd7058, -32'd6064},
{-32'd12792, 32'd3886, 32'd9499, -32'd2515},
{-32'd2923, -32'd2510, -32'd7748, 32'd7848},
{-32'd7702, -32'd7516, -32'd6511, 32'd5664},
{32'd11740, 32'd3713, 32'd4834, -32'd6445},
{-32'd2322, 32'd5267, -32'd7058, -32'd1735},
{32'd9381, -32'd3661, -32'd5650, 32'd87},
{-32'd6694, -32'd1340, -32'd7354, -32'd629},
{32'd10708, 32'd6446, -32'd9325, -32'd3328},
{32'd14629, 32'd8471, 32'd89, 32'd2802},
{32'd5724, 32'd2188, -32'd6043, -32'd5988},
{-32'd1576, -32'd12682, -32'd6503, -32'd9669},
{32'd3063, 32'd551, 32'd3620, 32'd4671},
{32'd6326, 32'd695, -32'd3784, 32'd6495},
{32'd5112, 32'd1225, -32'd7381, -32'd12832},
{-32'd6895, 32'd1748, -32'd2910, 32'd7210},
{32'd2743, 32'd4722, -32'd12958, 32'd938},
{-32'd4180, -32'd2629, 32'd2004, -32'd7204},
{32'd7407, 32'd1912, -32'd1419, -32'd5361},
{-32'd22301, -32'd4732, -32'd12599, -32'd3972},
{32'd647, 32'd6670, -32'd2223, -32'd9931},
{32'd1947, 32'd3237, -32'd10642, -32'd11100},
{32'd3321, -32'd32, -32'd464, 32'd1285},
{-32'd5387, -32'd8594, -32'd8605, -32'd1704},
{-32'd5241, -32'd2779, -32'd169, 32'd4919},
{32'd8303, 32'd1801, -32'd144, 32'd2956},
{-32'd7845, -32'd9986, -32'd2293, -32'd6280},
{32'd5826, -32'd7710, 32'd4581, -32'd2989},
{-32'd222, -32'd5667, 32'd7501, 32'd9178},
{-32'd804, 32'd11104, 32'd11446, 32'd571},
{-32'd2611, 32'd9779, -32'd3912, 32'd6784},
{32'd4869, 32'd3448, 32'd1722, -32'd6840},
{-32'd13656, -32'd5234, 32'd14305, -32'd1270},
{-32'd7261, 32'd5014, 32'd981, -32'd5766},
{-32'd4330, -32'd1736, -32'd4379, -32'd2404},
{-32'd2995, 32'd9078, -32'd7028, 32'd7893},
{32'd453, -32'd1609, -32'd421, 32'd1032},
{-32'd4294, 32'd6101, -32'd10346, -32'd8490},
{32'd2274, -32'd539, -32'd2085, 32'd2855},
{-32'd8661, 32'd593, 32'd7459, -32'd2290},
{-32'd2238, -32'd4005, 32'd2353, 32'd9179},
{32'd1061, -32'd4781, 32'd11186, 32'd449},
{32'd1539, -32'd7290, 32'd2054, -32'd6501},
{-32'd1694, 32'd5071, 32'd2312, 32'd2539},
{-32'd1987, 32'd3015, 32'd6797, 32'd1371},
{32'd4302, 32'd4627, -32'd9801, 32'd3712},
{-32'd12054, -32'd6341, -32'd1829, -32'd8630},
{32'd4360, 32'd294, -32'd923, -32'd2301},
{-32'd9508, -32'd7373, -32'd1621, -32'd5323},
{-32'd1380, -32'd6962, -32'd3989, 32'd1027},
{-32'd12512, 32'd9959, -32'd5126, -32'd4643},
{32'd8092, 32'd14042, 32'd10448, 32'd5061},
{32'd1932, -32'd5902, -32'd8329, 32'd7207},
{-32'd2921, -32'd8008, -32'd5999, -32'd1222},
{-32'd4089, -32'd5265, 32'd5242, -32'd3948},
{-32'd7406, 32'd786, 32'd2132, 32'd1588},
{-32'd2389, 32'd4970, 32'd10901, -32'd627},
{-32'd1125, -32'd1989, -32'd6341, -32'd1258},
{32'd4493, 32'd1805, 32'd14336, 32'd11890},
{32'd4191, -32'd3374, -32'd3977, 32'd2695},
{-32'd11929, 32'd6745, 32'd7498, 32'd573},
{32'd3750, 32'd2038, -32'd9584, 32'd3950},
{-32'd6780, 32'd7264, -32'd1474, -32'd2325},
{32'd3042, 32'd14705, -32'd12267, -32'd3400},
{32'd5160, 32'd2672, 32'd7656, 32'd11043},
{32'd109, -32'd600, -32'd4628, 32'd1004},
{32'd2, -32'd4219, -32'd7165, 32'd4350},
{-32'd4272, -32'd1489, 32'd4811, 32'd1322},
{32'd6392, -32'd12328, -32'd5135, -32'd13855},
{32'd3511, -32'd14184, -32'd5909, -32'd11209},
{32'd1518, 32'd8914, -32'd12264, -32'd7151},
{32'd9677, -32'd6165, 32'd1647, 32'd14007},
{-32'd5743, -32'd2581, 32'd15104, 32'd13253},
{-32'd316, 32'd2544, 32'd6842, 32'd1918},
{32'd481, 32'd2345, -32'd5740, -32'd14233},
{32'd4663, -32'd175, 32'd2333, -32'd8469},
{-32'd715, -32'd9213, -32'd9550, 32'd8922},
{-32'd2217, 32'd3990, 32'd4564, -32'd945},
{-32'd14624, -32'd2354, -32'd4803, 32'd7857},
{-32'd3999, 32'd5167, -32'd2580, 32'd6324},
{32'd1746, -32'd16812, -32'd9703, -32'd1568},
{-32'd4950, 32'd8062, 32'd4485, 32'd2471},
{-32'd6085, -32'd7175, -32'd4187, -32'd4249},
{32'd9969, 32'd6082, 32'd15140, 32'd7025},
{-32'd3102, -32'd8315, -32'd15268, -32'd3170},
{32'd2337, -32'd2069, -32'd10125, -32'd2706},
{32'd5463, 32'd4051, -32'd8970, -32'd5200},
{-32'd8878, -32'd5118, 32'd5737, 32'd362},
{-32'd16036, 32'd230, 32'd10531, -32'd8029},
{32'd1729, 32'd1023, 32'd9869, 32'd7799},
{-32'd5391, 32'd3575, -32'd261, -32'd4358},
{32'd9232, -32'd1219, 32'd2730, 32'd4497},
{32'd4276, 32'd5784, -32'd5775, -32'd2149},
{32'd8442, 32'd5574, -32'd2441, 32'd8033},
{-32'd8367, -32'd2033, -32'd11128, 32'd8120},
{32'd2104, -32'd17367, -32'd278, -32'd5977},
{32'd6209, 32'd6731, -32'd3330, -32'd4169},
{32'd7145, -32'd1969, 32'd5446, 32'd2042},
{32'd3612, 32'd9898, 32'd11911, 32'd6072},
{-32'd1561, 32'd4445, -32'd4870, 32'd1066},
{32'd1979, -32'd3207, -32'd2966, -32'd12978},
{32'd5129, -32'd7769, -32'd1189, -32'd3463},
{-32'd14569, -32'd7454, 32'd6248, -32'd32},
{32'd8153, 32'd2115, 32'd658, -32'd6877},
{32'd5735, 32'd969, 32'd1755, -32'd1641},
{32'd8277, 32'd10459, 32'd8200, 32'd8650},
{32'd8039, 32'd4856, 32'd855, 32'd1358}
},
{{-32'd125, 32'd5662, 32'd10746, -32'd2875},
{-32'd11383, -32'd7522, -32'd14893, -32'd5636},
{32'd1859, -32'd5218, -32'd10368, -32'd6726},
{32'd4305, 32'd7931, 32'd251, -32'd3720},
{-32'd3201, -32'd3257, 32'd2340, -32'd3965},
{32'd3948, -32'd11928, 32'd926, 32'd5154},
{-32'd379, 32'd2180, 32'd3924, 32'd5688},
{-32'd1253, 32'd1559, -32'd6654, -32'd1652},
{-32'd4778, -32'd2992, 32'd8605, -32'd1635},
{32'd8251, 32'd3811, 32'd5192, 32'd2861},
{-32'd8666, -32'd3610, 32'd183, -32'd1234},
{32'd3787, -32'd1987, -32'd4525, 32'd6862},
{-32'd2516, -32'd1403, 32'd7069, -32'd3252},
{-32'd2869, -32'd8530, -32'd6315, -32'd44},
{-32'd11225, 32'd5388, -32'd5902, -32'd5507},
{-32'd6883, 32'd4829, 32'd10832, -32'd7268},
{32'd10195, 32'd1463, 32'd6304, 32'd4594},
{-32'd5965, -32'd1824, 32'd1299, -32'd9020},
{32'd440, -32'd3713, 32'd272, -32'd8388},
{32'd6079, -32'd7686, -32'd4529, -32'd1688},
{32'd6526, 32'd5206, 32'd5244, -32'd15},
{-32'd1259, -32'd4091, -32'd2272, -32'd2035},
{-32'd4090, -32'd1251, 32'd725, -32'd1716},
{-32'd11124, -32'd478, -32'd1620, -32'd6651},
{32'd1591, -32'd2441, 32'd1849, -32'd859},
{32'd7016, -32'd4792, -32'd2100, -32'd3739},
{32'd198, -32'd6551, -32'd2312, 32'd496},
{-32'd444, 32'd2527, -32'd1309, -32'd4765},
{32'd622, 32'd1362, -32'd3, 32'd327},
{-32'd774, 32'd44, -32'd4215, 32'd1459},
{-32'd4292, -32'd7450, 32'd4342, -32'd2647},
{-32'd3306, -32'd9619, -32'd1841, -32'd3215},
{-32'd832, 32'd1503, -32'd1013, 32'd5027},
{-32'd3689, 32'd3491, -32'd754, -32'd3219},
{32'd5225, 32'd5978, 32'd5388, 32'd6702},
{-32'd2004, -32'd1578, 32'd5874, -32'd3601},
{32'd1494, -32'd4820, -32'd1367, -32'd4763},
{-32'd1205, -32'd4601, -32'd6253, 32'd4319},
{-32'd493, 32'd2882, -32'd39, 32'd879},
{-32'd283, 32'd10118, 32'd161, 32'd4145},
{32'd4983, 32'd3520, 32'd6165, 32'd10652},
{32'd3212, 32'd5084, 32'd8691, -32'd2225},
{-32'd9956, -32'd2486, 32'd3100, -32'd5379},
{-32'd7780, -32'd1016, -32'd592, -32'd8776},
{-32'd7582, -32'd2014, -32'd2648, -32'd642},
{32'd5580, -32'd4003, -32'd2184, 32'd601},
{-32'd7052, -32'd9205, -32'd9682, -32'd13740},
{-32'd1669, -32'd1110, -32'd4168, -32'd5504},
{32'd208, -32'd7122, 32'd7041, 32'd10352},
{32'd6172, -32'd3145, -32'd17482, -32'd4091},
{32'd4278, -32'd9568, -32'd63, 32'd2967},
{-32'd2947, 32'd1150, -32'd436, -32'd2171},
{-32'd4224, 32'd276, -32'd4357, -32'd10757},
{32'd912, 32'd2570, -32'd1604, -32'd706},
{-32'd2440, 32'd6337, 32'd6968, -32'd2016},
{-32'd1990, -32'd6091, -32'd4927, -32'd2160},
{32'd7854, 32'd3707, -32'd5021, 32'd5836},
{-32'd5417, -32'd13803, -32'd1858, -32'd5702},
{-32'd7984, 32'd2498, -32'd9780, -32'd773},
{32'd1639, -32'd1348, 32'd2409, 32'd6327},
{-32'd5345, 32'd1649, -32'd1168, 32'd906},
{-32'd5175, 32'd1673, -32'd7187, 32'd1034},
{-32'd11385, -32'd8029, 32'd1126, -32'd8130},
{32'd1082, -32'd7269, -32'd232, -32'd3163},
{-32'd5164, 32'd3336, -32'd2739, -32'd4714},
{32'd8013, 32'd1506, 32'd3679, -32'd388},
{32'd4725, -32'd364, -32'd3117, 32'd2324},
{32'd198, -32'd1340, -32'd13399, -32'd2077},
{-32'd377, 32'd11327, -32'd2381, -32'd8879},
{32'd8289, 32'd9597, -32'd6988, 32'd11645},
{32'd3581, -32'd700, 32'd1829, 32'd6978},
{-32'd66, -32'd1128, 32'd266, -32'd7664},
{-32'd5544, -32'd4163, 32'd3250, -32'd6467},
{32'd954, -32'd1391, 32'd1776, 32'd4233},
{32'd6363, 32'd6382, 32'd4722, 32'd17318},
{-32'd5389, 32'd13347, -32'd2161, -32'd7620},
{-32'd13274, -32'd1560, -32'd12119, -32'd3944},
{-32'd4517, -32'd1249, 32'd7131, -32'd1821},
{32'd635, 32'd5993, 32'd8735, 32'd13},
{-32'd2790, 32'd5319, 32'd4095, -32'd787},
{32'd455, 32'd3815, -32'd1728, 32'd1896},
{32'd5367, -32'd4515, 32'd17649, -32'd2288},
{32'd1070, -32'd3993, 32'd3663, -32'd2440},
{-32'd4249, 32'd522, -32'd253, -32'd6138},
{-32'd3732, 32'd4649, 32'd1709, -32'd10831},
{-32'd1648, -32'd6455, 32'd7443, -32'd375},
{-32'd1705, 32'd1497, 32'd1090, -32'd6910},
{-32'd8398, -32'd3470, 32'd8403, 32'd2424},
{32'd368, -32'd4248, -32'd2762, -32'd7664},
{32'd86, 32'd2571, -32'd1844, -32'd6639},
{32'd2948, 32'd1857, -32'd4869, 32'd2483},
{-32'd3223, -32'd2463, -32'd5093, -32'd5682},
{-32'd1451, 32'd1096, -32'd1454, -32'd4286},
{-32'd1841, 32'd4820, 32'd2107, 32'd2061},
{-32'd10017, -32'd7944, -32'd1657, -32'd5470},
{-32'd8012, -32'd762, -32'd10449, -32'd4179},
{32'd999, 32'd7107, 32'd4839, 32'd1140},
{32'd5693, 32'd6715, 32'd4986, 32'd3928},
{-32'd1707, -32'd828, 32'd10696, -32'd1850},
{32'd6896, 32'd4160, 32'd6317, 32'd4375},
{32'd1815, -32'd3394, -32'd6503, -32'd1882},
{-32'd162, -32'd1738, 32'd2940, -32'd2559},
{-32'd347, 32'd915, -32'd4907, 32'd2569},
{32'd7114, 32'd9683, 32'd8907, 32'd5442},
{32'd3758, -32'd2439, -32'd3169, 32'd1801},
{-32'd9664, -32'd1300, 32'd4770, -32'd7723},
{32'd764, -32'd9465, -32'd6289, 32'd9108},
{-32'd3759, 32'd1230, -32'd7718, 32'd6268},
{32'd10637, 32'd331, 32'd5022, 32'd7747},
{-32'd4228, -32'd163, -32'd9753, 32'd373},
{-32'd4248, 32'd9393, 32'd126, -32'd229},
{-32'd582, 32'd3114, 32'd7071, -32'd1674},
{-32'd1418, 32'd2275, 32'd526, 32'd1308},
{32'd3092, 32'd7399, 32'd5401, 32'd2154},
{-32'd7520, 32'd1873, 32'd613, -32'd4840},
{32'd2284, -32'd3903, -32'd453, 32'd1235},
{32'd6817, 32'd2287, 32'd211, 32'd3292},
{-32'd1314, 32'd9629, -32'd8554, -32'd1264},
{-32'd770, 32'd1023, 32'd7540, -32'd2979},
{32'd3249, 32'd4657, 32'd2974, 32'd2734},
{32'd5763, 32'd7315, 32'd3190, -32'd9359},
{32'd2631, 32'd4043, -32'd4419, -32'd5225},
{32'd10034, 32'd7441, -32'd6682, 32'd508},
{-32'd1954, -32'd2854, -32'd2473, -32'd977},
{-32'd1732, -32'd7698, 32'd820, -32'd4036},
{-32'd1607, -32'd6401, -32'd5788, 32'd7121},
{-32'd3393, 32'd1442, 32'd2357, 32'd4025},
{-32'd1458, -32'd4926, -32'd2104, -32'd2821},
{-32'd14522, -32'd1392, -32'd6309, 32'd2800},
{-32'd1443, -32'd13, 32'd2603, -32'd526},
{32'd3389, 32'd2433, 32'd7321, -32'd223},
{32'd967, -32'd2483, -32'd7973, 32'd7165},
{-32'd2587, -32'd4482, -32'd5741, -32'd5465},
{32'd1555, -32'd9991, -32'd3091, 32'd7811},
{32'd975, 32'd3858, 32'd3067, 32'd4093},
{-32'd982, 32'd2412, 32'd5811, -32'd245},
{-32'd10634, 32'd3574, 32'd8682, -32'd453},
{32'd1403, -32'd1786, -32'd5582, -32'd13046},
{32'd3414, 32'd1653, 32'd5088, 32'd7315},
{-32'd4768, -32'd1621, -32'd7287, -32'd2335},
{-32'd2349, 32'd613, -32'd1948, 32'd6150},
{-32'd1485, -32'd3579, -32'd215, -32'd3108},
{-32'd1115, 32'd2207, -32'd743, -32'd5847},
{32'd3009, -32'd6066, 32'd6470, -32'd1260},
{-32'd1833, 32'd3488, 32'd2993, -32'd1761},
{-32'd938, 32'd1835, -32'd2814, -32'd592},
{-32'd1921, -32'd3900, -32'd6411, 32'd4267},
{32'd6243, -32'd6442, 32'd2126, 32'd24},
{32'd5304, 32'd8914, 32'd4529, 32'd4918},
{-32'd2762, -32'd6140, -32'd5558, -32'd3699},
{-32'd9471, -32'd1874, -32'd327, -32'd8824},
{-32'd7609, 32'd3335, -32'd690, 32'd3527},
{32'd5397, 32'd1390, 32'd12045, -32'd13406},
{32'd6800, -32'd3455, -32'd2534, -32'd2866},
{-32'd2297, -32'd11147, -32'd2214, -32'd2485},
{-32'd8797, 32'd6881, 32'd5804, -32'd3584},
{-32'd30, 32'd5642, 32'd7447, 32'd5928},
{-32'd1601, 32'd993, -32'd5962, 32'd2454},
{-32'd613, -32'd3268, 32'd3664, 32'd1389},
{32'd408, 32'd1437, 32'd2449, -32'd751},
{32'd428, 32'd3693, -32'd3530, -32'd8731},
{-32'd3015, 32'd628, 32'd1108, -32'd7608},
{-32'd2971, -32'd611, 32'd736, -32'd2079},
{32'd1586, 32'd6967, -32'd5631, 32'd10953},
{-32'd90, 32'd2666, -32'd4025, 32'd8711},
{32'd757, -32'd4484, -32'd2630, 32'd1975},
{-32'd2602, -32'd14583, 32'd34, -32'd2461},
{-32'd10684, -32'd4456, -32'd4364, 32'd697},
{-32'd4989, 32'd5115, -32'd1403, -32'd7983},
{-32'd5846, 32'd374, -32'd2246, -32'd247},
{-32'd6259, -32'd2482, 32'd1124, 32'd2205},
{32'd3127, -32'd244, -32'd7175, 32'd10742},
{32'd7367, 32'd9093, 32'd2903, 32'd7850},
{-32'd706, -32'd1885, -32'd2016, 32'd2209},
{32'd9753, -32'd5367, 32'd5850, -32'd1130},
{32'd3292, -32'd5052, 32'd6182, -32'd1124},
{32'd2523, 32'd4955, -32'd5444, 32'd15916},
{32'd4632, -32'd359, -32'd8577, 32'd9307},
{-32'd8694, 32'd5961, 32'd6450, 32'd1017},
{-32'd3618, -32'd5214, -32'd9974, 32'd1234},
{-32'd3867, 32'd5128, -32'd2539, -32'd7675},
{-32'd7494, -32'd1958, -32'd3381, -32'd4867},
{32'd545, -32'd1154, -32'd356, -32'd10222},
{-32'd504, -32'd6990, 32'd595, -32'd918},
{-32'd8832, -32'd6078, -32'd15341, -32'd1561},
{32'd12585, -32'd2572, -32'd1187, 32'd11976},
{-32'd650, 32'd9207, -32'd1230, 32'd4256},
{32'd9176, 32'd5535, 32'd1386, 32'd3382},
{-32'd2619, -32'd6034, 32'd1324, 32'd7527},
{32'd6081, -32'd4280, 32'd3938, -32'd1182},
{-32'd1228, 32'd1097, 32'd1084, -32'd2860},
{-32'd13889, -32'd8199, -32'd3044, -32'd501},
{32'd951, -32'd4136, -32'd6159, 32'd5362},
{32'd5640, -32'd4675, 32'd6408, -32'd4115},
{32'd9645, -32'd94, -32'd1765, -32'd2359},
{-32'd1260, -32'd6040, 32'd5886, 32'd1287},
{-32'd1625, 32'd900, -32'd714, 32'd10963},
{32'd2846, 32'd1801, 32'd6466, 32'd1036},
{-32'd2637, 32'd1486, -32'd4957, 32'd15142},
{-32'd256, 32'd2950, -32'd4926, -32'd8190},
{-32'd5055, -32'd6749, -32'd9482, -32'd1818},
{-32'd6188, 32'd1262, -32'd483, 32'd3504},
{32'd1411, -32'd5721, 32'd5882, 32'd14231},
{-32'd8773, 32'd3410, 32'd4707, 32'd4584},
{-32'd5839, -32'd5345, -32'd1894, -32'd9910},
{-32'd4046, -32'd5022, -32'd7631, 32'd698},
{32'd2132, 32'd10177, 32'd3439, 32'd5344},
{-32'd4240, 32'd1754, -32'd554, -32'd9218},
{-32'd11900, 32'd2635, 32'd9806, -32'd7079},
{-32'd8, 32'd3684, -32'd185, -32'd4378},
{-32'd6287, 32'd1375, -32'd1130, -32'd4275},
{32'd3665, -32'd1229, -32'd2182, 32'd261},
{-32'd1929, -32'd847, -32'd7785, 32'd1010},
{32'd10711, 32'd2704, -32'd249, 32'd8693},
{-32'd5570, 32'd2505, -32'd8072, -32'd10664},
{-32'd1758, 32'd1293, 32'd2013, -32'd3136},
{32'd5563, 32'd545, 32'd2846, 32'd6209},
{32'd1356, -32'd6371, -32'd6000, -32'd4002},
{32'd4717, 32'd9185, 32'd3281, 32'd3786},
{-32'd1086, 32'd7174, 32'd286, -32'd7829},
{32'd4795, -32'd3985, -32'd560, 32'd1865},
{32'd197, 32'd3480, 32'd343, 32'd953},
{32'd7031, 32'd687, 32'd4606, 32'd3738},
{32'd5031, -32'd618, 32'd9819, 32'd2372},
{32'd4389, -32'd1217, -32'd801, -32'd1845},
{32'd2767, 32'd4879, 32'd2597, 32'd7870},
{-32'd5100, 32'd5528, -32'd1016, 32'd2922},
{-32'd3076, -32'd1590, -32'd961, -32'd7873},
{32'd1387, 32'd12789, 32'd1289, -32'd7649},
{32'd4195, 32'd3803, -32'd3056, -32'd7096},
{32'd6726, 32'd5807, -32'd5517, 32'd3397},
{32'd2373, -32'd5153, -32'd839, -32'd562},
{-32'd120, 32'd6128, 32'd4340, 32'd1222},
{-32'd6233, 32'd3003, -32'd2160, -32'd12863},
{-32'd3965, -32'd8688, -32'd5750, -32'd6811},
{-32'd8101, -32'd14312, -32'd7459, -32'd3630},
{32'd623, 32'd3397, -32'd7460, -32'd780},
{32'd5491, -32'd3712, -32'd872, 32'd6504},
{32'd9840, 32'd3453, 32'd3158, 32'd13036},
{-32'd8315, -32'd5649, -32'd3568, -32'd9031},
{-32'd2061, -32'd3804, 32'd997, -32'd2463},
{-32'd5965, -32'd1848, -32'd846, -32'd15422},
{-32'd12665, -32'd4552, -32'd5896, -32'd5130},
{-32'd9460, -32'd3843, -32'd4644, 32'd6130},
{32'd8792, 32'd11187, 32'd5587, 32'd5377},
{-32'd5837, 32'd5038, 32'd7389, 32'd6136},
{-32'd6274, -32'd529, -32'd2516, -32'd6730},
{32'd8161, -32'd12033, -32'd3801, 32'd5260},
{32'd6180, 32'd2188, 32'd6433, -32'd5434},
{-32'd9305, -32'd6215, 32'd2918, 32'd2318},
{-32'd6562, -32'd5154, 32'd1629, -32'd14934},
{-32'd2619, 32'd2139, -32'd4415, 32'd4099},
{-32'd537, -32'd1148, -32'd357, 32'd4378},
{32'd389, -32'd362, -32'd5063, -32'd768},
{-32'd57, 32'd695, -32'd1038, 32'd4155},
{-32'd3814, 32'd1060, 32'd3741, 32'd10230},
{-32'd1391, -32'd16137, -32'd78, 32'd8821},
{32'd7967, 32'd7181, -32'd597, -32'd1731},
{-32'd7229, -32'd142, 32'd2408, -32'd3525},
{32'd6611, -32'd7708, 32'd6123, 32'd5861},
{32'd4499, -32'd9119, 32'd5918, 32'd12922},
{-32'd1429, 32'd3957, 32'd5946, 32'd1832},
{-32'd537, -32'd5543, -32'd6178, -32'd9610},
{-32'd733, 32'd1880, -32'd11382, -32'd3124},
{32'd5586, 32'd6335, -32'd2844, -32'd3205},
{32'd5413, -32'd5263, -32'd5102, 32'd491},
{32'd4244, -32'd123, 32'd667, 32'd3962},
{-32'd6418, 32'd3669, -32'd276, -32'd10533},
{-32'd7026, -32'd6852, -32'd2770, 32'd1567},
{-32'd11072, -32'd9405, -32'd4583, -32'd511},
{32'd427, 32'd10592, 32'd6618, -32'd1500},
{32'd9122, -32'd253, -32'd1339, -32'd903},
{32'd5865, -32'd9835, -32'd1083, 32'd6905},
{-32'd1628, -32'd3130, 32'd868, -32'd354},
{-32'd1133, -32'd3862, -32'd4535, -32'd2976},
{-32'd8879, -32'd5118, 32'd3719, 32'd968},
{32'd6959, 32'd5950, 32'd5711, 32'd3190},
{-32'd2073, 32'd4496, 32'd4726, -32'd3459},
{-32'd4352, -32'd1806, 32'd1488, -32'd859},
{-32'd656, 32'd2009, -32'd4779, -32'd3271},
{32'd5279, 32'd906, 32'd1803, 32'd4485},
{32'd1561, -32'd5224, -32'd7609, 32'd23869},
{32'd1063, -32'd3568, 32'd7432, 32'd5920},
{32'd333, -32'd5901, -32'd3173, 32'd4617},
{32'd8790, 32'd1191, 32'd6615, -32'd885},
{-32'd1941, -32'd1797, -32'd11685, -32'd11688},
{32'd6408, -32'd10627, 32'd3078, 32'd5579},
{-32'd611, -32'd2870, -32'd4750, -32'd6038},
{-32'd1500, 32'd3910, 32'd1949, -32'd13457},
{-32'd7833, 32'd4901, -32'd9778, 32'd5889},
{32'd263, -32'd406, 32'd11599, -32'd3807},
{32'd5003, 32'd6401, 32'd2203, 32'd2805},
{32'd629, 32'd2847, 32'd2980, 32'd2494},
{32'd3922, 32'd2719, -32'd2249, 32'd1481},
{-32'd289, -32'd3090, -32'd419, 32'd3931},
{-32'd793, 32'd3688, -32'd4300, -32'd2588},
{-32'd4224, -32'd3807, -32'd3867, 32'd5057},
{-32'd2833, 32'd6368, 32'd6616, -32'd1770},
{32'd3717, 32'd10100, 32'd6273, 32'd4093},
{-32'd6724, -32'd5129, -32'd1102, 32'd1169}
},
{{32'd12418, 32'd4204, 32'd968, -32'd920},
{-32'd2900, 32'd1987, -32'd2569, -32'd1865},
{-32'd1640, -32'd3395, -32'd807, -32'd1561},
{32'd7250, 32'd5804, 32'd5016, 32'd6831},
{-32'd1977, -32'd5760, 32'd604, -32'd7685},
{-32'd196, -32'd305, -32'd323, 32'd7301},
{-32'd764, -32'd8472, 32'd3348, 32'd921},
{32'd5129, -32'd997, -32'd2899, -32'd4420},
{-32'd11377, 32'd2634, 32'd2485, 32'd1056},
{32'd8549, 32'd6722, 32'd5043, 32'd2952},
{-32'd15561, -32'd10399, 32'd697, 32'd7606},
{32'd11660, 32'd4392, 32'd5650, 32'd12613},
{32'd7095, 32'd424, -32'd296, -32'd3620},
{-32'd5646, -32'd5484, -32'd12049, -32'd1142},
{32'd5438, -32'd1731, 32'd110, 32'd7725},
{-32'd6717, -32'd5001, -32'd4285, -32'd5957},
{32'd7841, 32'd7007, -32'd1206, 32'd2087},
{32'd5344, 32'd2937, -32'd720, 32'd1292},
{-32'd4099, -32'd2443, -32'd4638, 32'd1833},
{32'd1580, 32'd1786, -32'd9745, -32'd6183},
{-32'd5021, -32'd2233, 32'd3660, 32'd610},
{-32'd2749, 32'd3719, -32'd3935, -32'd8543},
{-32'd430, 32'd2994, -32'd4601, -32'd7974},
{-32'd7407, -32'd1768, -32'd5, 32'd2956},
{32'd8361, -32'd2210, 32'd9299, 32'd3885},
{32'd1253, 32'd13128, 32'd1063, 32'd3997},
{32'd3908, 32'd8235, 32'd9323, 32'd1243},
{32'd3902, -32'd1564, -32'd3280, 32'd3886},
{32'd9110, 32'd520, -32'd3403, 32'd11253},
{32'd4527, -32'd7870, -32'd7766, 32'd7889},
{32'd4308, -32'd8738, 32'd2873, 32'd2419},
{-32'd1417, -32'd7522, -32'd5621, 32'd408},
{-32'd1767, -32'd3487, -32'd805, 32'd2449},
{-32'd10588, -32'd2807, -32'd1848, -32'd1817},
{32'd10976, 32'd4823, 32'd7043, 32'd1766},
{-32'd10929, -32'd1848, -32'd6796, -32'd480},
{32'd5102, 32'd7863, -32'd3094, -32'd8996},
{32'd2453, 32'd627, -32'd17283, 32'd987},
{32'd8072, 32'd5029, 32'd2801, 32'd1128},
{32'd2536, 32'd2642, 32'd9154, -32'd746},
{-32'd1554, -32'd3423, -32'd3, -32'd4927},
{32'd5166, -32'd1680, 32'd2291, 32'd7524},
{-32'd4703, 32'd4012, -32'd518, -32'd3266},
{-32'd5292, -32'd8449, 32'd3238, -32'd6890},
{-32'd3536, -32'd3928, -32'd4905, -32'd9992},
{-32'd13096, 32'd4138, -32'd7672, -32'd2159},
{32'd522, -32'd9394, -32'd5853, -32'd7416},
{32'd5762, 32'd3226, -32'd5901, -32'd2786},
{32'd3320, 32'd3581, 32'd4165, 32'd7205},
{32'd2232, 32'd2053, -32'd1687, -32'd2548},
{-32'd3094, -32'd1876, 32'd1535, 32'd3157},
{32'd2994, 32'd4755, 32'd7883, 32'd4164},
{32'd3362, 32'd2119, 32'd7087, -32'd41},
{-32'd6863, -32'd17517, -32'd10079, -32'd7646},
{-32'd3230, -32'd1396, -32'd3361, -32'd5316},
{-32'd4318, 32'd763, -32'd3752, 32'd900},
{32'd223, -32'd1404, 32'd8493, -32'd1370},
{-32'd7777, -32'd10755, -32'd5449, -32'd1793},
{-32'd18549, 32'd4885, -32'd960, -32'd2014},
{32'd4620, 32'd6730, -32'd1844, 32'd1742},
{32'd4880, 32'd6685, -32'd2272, 32'd1049},
{-32'd10816, -32'd5426, 32'd173, -32'd982},
{32'd129, -32'd9347, -32'd4013, 32'd1677},
{32'd2956, 32'd1369, -32'd1484, -32'd5592},
{32'd1179, 32'd4101, 32'd8683, -32'd3489},
{32'd7904, 32'd1157, 32'd7331, 32'd2776},
{32'd11510, 32'd16296, 32'd1209, -32'd803},
{32'd1862, 32'd3198, 32'd3272, 32'd2178},
{32'd12042, -32'd1047, -32'd4738, 32'd6879},
{32'd3418, -32'd917, 32'd1273, 32'd12194},
{-32'd66, -32'd44, 32'd1321, -32'd9810},
{32'd1305, -32'd10302, -32'd5400, 32'd3671},
{-32'd12814, -32'd7792, -32'd2654, -32'd2356},
{-32'd3134, -32'd3821, 32'd3412, -32'd553},
{32'd6725, 32'd8243, 32'd2184, 32'd5754},
{32'd1537, -32'd5515, -32'd5628, -32'd15433},
{-32'd4658, -32'd10142, 32'd2652, -32'd1592},
{-32'd2004, 32'd13821, -32'd2813, 32'd8819},
{32'd9469, 32'd3574, 32'd11970, 32'd5631},
{-32'd3355, -32'd6977, -32'd5550, -32'd475},
{32'd10913, 32'd3211, 32'd6122, -32'd3271},
{32'd4293, 32'd4016, -32'd2806, -32'd5832},
{-32'd7048, -32'd2589, 32'd4369, -32'd6581},
{32'd4075, -32'd714, 32'd13414, -32'd6418},
{32'd9451, -32'd8522, -32'd7619, -32'd9578},
{32'd2150, 32'd763, -32'd7674, -32'd3086},
{32'd3315, 32'd4711, -32'd15104, -32'd3625},
{-32'd12207, -32'd12514, -32'd17065, -32'd10029},
{32'd1394, -32'd4131, -32'd4314, 32'd8348},
{32'd1631, 32'd59, 32'd113, -32'd4100},
{32'd2897, -32'd4965, 32'd3091, 32'd1659},
{-32'd494, -32'd390, 32'd3155, -32'd3058},
{32'd10118, -32'd3418, -32'd3353, 32'd3456},
{32'd4153, 32'd18105, 32'd2511, -32'd357},
{32'd1638, 32'd889, 32'd2455, -32'd277},
{-32'd280, -32'd5493, 32'd2395, -32'd13016},
{32'd8754, 32'd2366, -32'd2351, 32'd5761},
{-32'd81, 32'd298, 32'd5060, -32'd1061},
{-32'd3506, -32'd749, -32'd2817, 32'd908},
{32'd14139, 32'd6091, 32'd4121, 32'd164},
{32'd5493, -32'd1295, -32'd9684, 32'd4484},
{-32'd481, -32'd3098, 32'd1773, -32'd10436},
{32'd1698, -32'd8216, 32'd373, -32'd2275},
{32'd768, 32'd558, 32'd1235, 32'd1447},
{-32'd4485, -32'd152, 32'd4468, 32'd6560},
{32'd4669, 32'd2075, 32'd3434, 32'd3507},
{-32'd17803, -32'd4487, 32'd2153, 32'd8625},
{-32'd1416, -32'd2034, 32'd17492, -32'd7491},
{32'd7692, 32'd13643, 32'd2961, -32'd573},
{-32'd5450, 32'd70, -32'd2237, -32'd13891},
{-32'd8403, -32'd676, 32'd8968, -32'd1273},
{32'd6234, -32'd373, -32'd4138, -32'd1975},
{32'd5695, 32'd5403, 32'd5850, -32'd6567},
{32'd1782, 32'd3806, -32'd1820, -32'd11354},
{-32'd11467, 32'd230, -32'd7904, -32'd1508},
{-32'd8230, 32'd1638, 32'd3124, -32'd5998},
{32'd947, 32'd1093, 32'd13313, 32'd8373},
{32'd3922, -32'd2776, 32'd7053, 32'd3532},
{-32'd6743, -32'd11213, 32'd1301, 32'd7466},
{32'd7483, 32'd9303, 32'd12330, 32'd9338},
{-32'd2615, 32'd3515, 32'd1719, -32'd11588},
{-32'd253, -32'd3091, 32'd10833, 32'd3745},
{32'd225, -32'd600, 32'd264, 32'd671},
{32'd3175, 32'd1890, -32'd6838, -32'd3353},
{32'd6666, -32'd3848, -32'd5984, -32'd4422},
{32'd6189, 32'd4383, 32'd11525, -32'd149},
{-32'd2587, -32'd745, -32'd6939, -32'd7000},
{-32'd1470, 32'd177, 32'd1969, -32'd3711},
{-32'd3734, 32'd9388, -32'd2141, 32'd645},
{-32'd7340, -32'd2100, 32'd6528, 32'd1707},
{32'd494, -32'd7454, -32'd6184, -32'd5836},
{32'd2464, -32'd15705, -32'd5960, 32'd1982},
{-32'd869, -32'd3221, 32'd1216, 32'd3299},
{-32'd200, -32'd3543, 32'd7517, -32'd8073},
{32'd8960, -32'd2111, -32'd2596, 32'd1966},
{-32'd1249, 32'd4106, -32'd1059, -32'd4676},
{32'd1696, -32'd6865, -32'd8719, 32'd942},
{-32'd5277, 32'd2002, 32'd1965, -32'd1052},
{32'd11178, 32'd246, -32'd113, 32'd6373},
{-32'd3610, -32'd1215, -32'd7932, -32'd8167},
{-32'd8692, 32'd3263, -32'd768, 32'd2399},
{-32'd585, -32'd6788, -32'd4348, -32'd10474},
{-32'd2166, 32'd910, -32'd1955, 32'd3731},
{-32'd793, -32'd2369, -32'd13519, -32'd3267},
{32'd11368, 32'd9402, 32'd3385, -32'd4476},
{32'd6677, 32'd2816, 32'd5374, -32'd4216},
{-32'd3279, -32'd10345, -32'd5585, -32'd6586},
{-32'd3814, -32'd3160, -32'd611, -32'd1405},
{32'd5770, -32'd1326, 32'd4148, 32'd2826},
{-32'd2718, -32'd6262, -32'd3238, -32'd4530},
{-32'd11203, -32'd5965, -32'd3663, 32'd2227},
{32'd7159, -32'd1154, -32'd4089, -32'd5055},
{32'd1805, -32'd3189, 32'd522, -32'd3353},
{32'd2929, 32'd1317, -32'd3154, -32'd18988},
{-32'd6670, -32'd7948, 32'd1674, -32'd4021},
{32'd3711, -32'd4057, -32'd1080, 32'd2435},
{-32'd5595, 32'd5039, -32'd2696, 32'd2299},
{32'd1189, 32'd4200, 32'd5096, 32'd6181},
{32'd2580, -32'd4087, 32'd2844, 32'd4017},
{32'd777, -32'd3163, -32'd486, 32'd105},
{-32'd11415, -32'd6552, 32'd802, 32'd9},
{32'd2499, 32'd202, 32'd6537, -32'd2889},
{-32'd16235, -32'd5534, -32'd11678, -32'd6177},
{32'd5513, 32'd2834, 32'd5871, 32'd9483},
{32'd907, 32'd2136, 32'd1943, -32'd527},
{32'd5153, 32'd4875, 32'd8924, -32'd4270},
{-32'd441, -32'd4497, 32'd11308, -32'd2294},
{-32'd879, -32'd4049, -32'd5779, 32'd7226},
{-32'd8502, -32'd1032, -32'd8911, -32'd5395},
{-32'd8304, -32'd14496, -32'd9269, -32'd2761},
{-32'd5269, -32'd6032, 32'd11595, 32'd7750},
{-32'd2168, -32'd5760, 32'd8717, 32'd7736},
{32'd8153, 32'd7386, 32'd9738, -32'd445},
{-32'd10160, -32'd6099, -32'd11153, 32'd2821},
{32'd7896, 32'd960, 32'd4579, 32'd13288},
{32'd263, -32'd22, -32'd2638, -32'd12123},
{32'd2317, -32'd4046, -32'd316, -32'd10556},
{32'd4145, -32'd1815, -32'd3118, -32'd990},
{32'd3305, -32'd1492, -32'd5911, -32'd7887},
{-32'd716, 32'd236, -32'd5661, 32'd1833},
{-32'd6348, -32'd1564, -32'd7480, -32'd1684},
{-32'd12537, -32'd10014, -32'd4291, -32'd2663},
{-32'd1192, 32'd317, -32'd2199, 32'd4760},
{32'd6751, 32'd92, 32'd793, -32'd687},
{32'd1223, -32'd6440, 32'd1248, 32'd3925},
{32'd4039, 32'd8233, 32'd7874, 32'd2343},
{32'd12455, 32'd4430, 32'd8055, 32'd9461},
{-32'd4554, -32'd2867, 32'd6518, 32'd10372},
{32'd2150, -32'd1534, 32'd1086, 32'd988},
{-32'd14635, -32'd3418, -32'd59, 32'd5598},
{-32'd216, 32'd768, 32'd1218, -32'd3081},
{-32'd16209, -32'd10798, -32'd3105, 32'd1292},
{32'd9178, 32'd7265, 32'd8268, 32'd9277},
{-32'd675, 32'd3894, 32'd5908, 32'd99},
{32'd4136, -32'd9025, 32'd1023, -32'd4686},
{32'd5669, 32'd8124, -32'd9075, -32'd9771},
{32'd4149, 32'd3945, -32'd580, -32'd2760},
{-32'd7035, 32'd7008, 32'd3357, 32'd2598},
{-32'd8114, -32'd6511, 32'd1739, 32'd2000},
{-32'd4639, -32'd3289, 32'd8600, -32'd7459},
{-32'd10602, -32'd8780, -32'd12687, -32'd4384},
{32'd649, -32'd1609, 32'd4216, -32'd5890},
{32'd4290, 32'd714, -32'd2463, -32'd12411},
{32'd7885, 32'd770, -32'd4335, 32'd2610},
{32'd3773, 32'd4225, 32'd2211, 32'd6963},
{-32'd2451, 32'd11057, -32'd9010, 32'd7310},
{32'd4846, 32'd1120, 32'd7995, 32'd1191},
{-32'd173, 32'd24, -32'd2535, -32'd2310},
{32'd7287, 32'd4443, -32'd10775, 32'd1257},
{32'd154, 32'd730, 32'd2963, -32'd1419},
{-32'd6906, -32'd3108, 32'd7102, 32'd4388},
{-32'd4676, 32'd5921, 32'd986, -32'd6495},
{-32'd6344, -32'd12665, -32'd4130, -32'd9583},
{32'd3000, 32'd7077, 32'd1120, 32'd14420},
{-32'd11965, 32'd6364, -32'd6471, -32'd14569},
{32'd8707, -32'd2814, -32'd11052, 32'd3797},
{32'd12407, 32'd3001, 32'd822, -32'd1615},
{32'd4926, -32'd11543, 32'd9649, 32'd9701},
{-32'd1662, 32'd11898, -32'd1375, 32'd5692},
{32'd920, -32'd4199, 32'd6890, 32'd5676},
{-32'd5714, -32'd7946, -32'd4439, 32'd8846},
{-32'd932, -32'd3758, 32'd8369, 32'd8588},
{32'd1716, 32'd9191, 32'd12584, 32'd347},
{-32'd5632, -32'd6855, -32'd4710, 32'd326},
{-32'd872, -32'd3473, -32'd3207, -32'd4207},
{-32'd8591, -32'd2020, -32'd14722, -32'd5998},
{32'd5697, 32'd881, -32'd3685, 32'd8426},
{-32'd2455, 32'd6801, -32'd3710, 32'd1273},
{-32'd124, 32'd1579, -32'd2630, 32'd6047},
{-32'd725, 32'd1347, 32'd7815, 32'd7370},
{-32'd7031, -32'd11701, -32'd5307, 32'd7396},
{-32'd7943, -32'd10002, -32'd3782, -32'd4414},
{-32'd7257, -32'd7228, 32'd3911, 32'd13481},
{32'd1898, -32'd1344, -32'd1832, -32'd2391},
{-32'd3205, -32'd3475, -32'd4392, -32'd1071},
{-32'd6201, -32'd4939, -32'd5986, -32'd10659},
{-32'd3179, -32'd1345, -32'd6370, -32'd349},
{-32'd1783, -32'd7169, -32'd9438, 32'd5756},
{32'd4068, 32'd2681, 32'd7992, 32'd649},
{-32'd8313, 32'd316, 32'd3129, 32'd2236},
{-32'd2963, -32'd9429, -32'd2127, -32'd3189},
{-32'd4593, 32'd3546, -32'd2092, 32'd2170},
{-32'd9351, -32'd7136, -32'd401, -32'd5517},
{-32'd7544, 32'd2349, 32'd3512, 32'd4413},
{32'd3671, 32'd9581, 32'd7561, 32'd4577},
{32'd8869, -32'd510, -32'd3388, 32'd4450},
{32'd5925, -32'd6329, 32'd864, -32'd4673},
{32'd11740, -32'd162, -32'd1668, -32'd8909},
{-32'd1117, 32'd2756, 32'd1027, 32'd14270},
{-32'd8232, -32'd166, 32'd3628, 32'd142},
{-32'd1452, 32'd7494, -32'd738, -32'd3941},
{-32'd1136, 32'd5443, -32'd2137, 32'd1875},
{32'd6598, 32'd6735, 32'd42, 32'd2424},
{32'd2668, 32'd727, -32'd1656, 32'd287},
{-32'd9883, -32'd4915, -32'd15677, -32'd5377},
{32'd6358, 32'd4512, -32'd4861, -32'd4983},
{32'd22, 32'd5365, 32'd1623, -32'd9690},
{32'd19561, 32'd5369, -32'd2770, -32'd2940},
{-32'd16407, -32'd12441, -32'd10026, -32'd1502},
{-32'd3210, 32'd14076, -32'd249, 32'd72},
{32'd5019, 32'd564, -32'd767, 32'd678},
{32'd3220, 32'd4282, 32'd1188, -32'd6485},
{-32'd2684, -32'd1839, -32'd9605, 32'd6205},
{-32'd1964, 32'd3054, -32'd7353, -32'd1781},
{32'd4087, -32'd3045, 32'd16687, -32'd876},
{-32'd710, 32'd589, -32'd8673, 32'd212},
{-32'd2879, -32'd1811, 32'd3053, 32'd13546},
{-32'd6287, 32'd262, 32'd488, 32'd5051},
{-32'd1771, -32'd4427, -32'd6968, -32'd9230},
{-32'd10095, -32'd1377, -32'd5080, -32'd1465},
{32'd3093, 32'd2193, -32'd670, 32'd7989},
{32'd3036, -32'd162, 32'd3399, 32'd4266},
{32'd4360, 32'd437, -32'd6482, 32'd2591},
{-32'd16727, -32'd7806, 32'd6077, -32'd6422},
{32'd2819, 32'd1703, -32'd5497, 32'd2834},
{32'd2143, -32'd928, -32'd579, -32'd2170},
{32'd8120, 32'd8864, 32'd4762, 32'd4454},
{-32'd2930, 32'd2287, 32'd11163, 32'd4432},
{-32'd8499, -32'd2366, -32'd8053, 32'd910},
{32'd6475, -32'd98, 32'd1340, -32'd2543},
{32'd6751, -32'd1918, 32'd9366, 32'd848},
{-32'd4544, 32'd651, -32'd3699, -32'd8337},
{-32'd1349, 32'd3634, -32'd4239, -32'd2371},
{32'd3042, 32'd7708, 32'd5427, 32'd13639},
{32'd4335, 32'd9969, 32'd11774, -32'd5661},
{-32'd11647, -32'd3679, -32'd4145, -32'd5016},
{32'd5979, 32'd11570, 32'd1534, -32'd5417},
{-32'd3587, -32'd4865, -32'd5615, -32'd2121},
{32'd4078, 32'd7447, -32'd4486, 32'd1030},
{-32'd8912, -32'd7894, -32'd6350, 32'd563},
{-32'd2469, -32'd10025, 32'd1097, 32'd8656},
{-32'd3590, 32'd11464, 32'd5387, 32'd3085},
{-32'd4674, 32'd318, -32'd1545, -32'd12765},
{32'd826, -32'd5628, 32'd978, -32'd5237},
{-32'd1007, -32'd6724, -32'd4360, 32'd3586},
{-32'd5229, -32'd4338, -32'd3462, 32'd1073},
{-32'd4617, -32'd8660, 32'd3289, -32'd4626},
{32'd586, 32'd9977, 32'd972, -32'd931},
{32'd19746, 32'd4328, 32'd5288, -32'd1523},
{-32'd7529, -32'd11738, -32'd6823, -32'd4425}
},
{{32'd14368, -32'd4148, -32'd9262, -32'd1235},
{-32'd22245, -32'd15913, -32'd4260, 32'd4615},
{32'd5509, 32'd2082, 32'd2712, -32'd4408},
{-32'd4208, 32'd9312, 32'd1447, 32'd5953},
{-32'd3566, 32'd7460, 32'd9396, 32'd4971},
{-32'd5899, 32'd6273, 32'd4954, -32'd4410},
{-32'd2255, 32'd10617, 32'd1867, -32'd2413},
{-32'd191, 32'd9106, -32'd5027, 32'd9732},
{-32'd10059, 32'd10230, 32'd15522, 32'd5423},
{32'd8117, 32'd6551, -32'd169, 32'd2929},
{32'd1750, -32'd5727, -32'd8538, -32'd6517},
{32'd5168, -32'd5272, 32'd5197, 32'd1421},
{32'd1999, 32'd2702, -32'd11769, 32'd7556},
{-32'd2187, 32'd6596, 32'd5496, -32'd2212},
{-32'd3377, 32'd10796, -32'd11889, -32'd8149},
{32'd235, -32'd6907, -32'd11558, 32'd5854},
{-32'd6309, -32'd177, 32'd7812, 32'd7954},
{32'd7044, 32'd6631, -32'd6808, 32'd5565},
{-32'd8713, 32'd14740, -32'd14426, -32'd6868},
{-32'd824, 32'd3657, -32'd1316, 32'd7785},
{-32'd8960, -32'd7477, -32'd6506, -32'd2731},
{-32'd11031, 32'd1051, -32'd9224, -32'd10169},
{-32'd6671, 32'd6799, 32'd483, -32'd3726},
{32'd816, -32'd3219, -32'd12039, -32'd16585},
{32'd8920, 32'd2979, 32'd1844, -32'd7786},
{32'd6943, -32'd5392, 32'd8148, -32'd6225},
{-32'd1412, -32'd9648, -32'd15638, 32'd676},
{-32'd7444, 32'd8289, 32'd10632, 32'd2609},
{-32'd2765, 32'd6058, 32'd5315, -32'd6610},
{32'd3680, 32'd13360, 32'd9203, 32'd16434},
{32'd373, -32'd1980, 32'd890, 32'd7770},
{-32'd7417, 32'd3758, 32'd7232, -32'd9711},
{32'd8235, -32'd6564, 32'd2383, 32'd7853},
{32'd330, -32'd6277, -32'd2800, 32'd2546},
{32'd10613, 32'd11149, -32'd3105, -32'd2861},
{-32'd5875, -32'd7695, -32'd6700, 32'd7238},
{-32'd247, 32'd4383, 32'd12991, 32'd15780},
{-32'd1293, -32'd7321, 32'd10359, -32'd4312},
{-32'd10921, 32'd3932, 32'd5690, -32'd10617},
{32'd13099, 32'd7626, 32'd2347, 32'd10406},
{-32'd3678, -32'd6722, -32'd4193, -32'd11533},
{32'd801, 32'd2991, -32'd11555, 32'd8054},
{32'd4342, -32'd1740, 32'd776, -32'd3517},
{-32'd5926, -32'd3318, -32'd16084, 32'd1122},
{32'd4713, 32'd5128, -32'd3490, -32'd546},
{32'd14560, 32'd3551, 32'd10335, -32'd961},
{32'd650, 32'd9692, -32'd1466, 32'd9375},
{-32'd3614, -32'd8661, 32'd396, 32'd3014},
{32'd1003, 32'd9920, -32'd8035, -32'd13188},
{32'd2019, -32'd758, 32'd11336, -32'd4749},
{-32'd9767, -32'd9102, 32'd304, 32'd2009},
{32'd722, 32'd6548, -32'd9917, -32'd12057},
{32'd3847, -32'd2668, -32'd1559, -32'd2070},
{32'd2898, 32'd3490, -32'd1487, -32'd689},
{32'd292, 32'd2908, -32'd2901, -32'd2181},
{32'd958, -32'd8911, 32'd5620, 32'd13288},
{32'd7708, 32'd11508, 32'd5545, -32'd4162},
{32'd7773, -32'd5250, 32'd2166, -32'd8830},
{-32'd5570, 32'd3980, -32'd4605, -32'd4927},
{32'd8014, 32'd808, -32'd5020, 32'd7632},
{-32'd3094, 32'd105, -32'd2053, 32'd7077},
{32'd4217, 32'd3198, 32'd18343, 32'd14135},
{-32'd264, -32'd3285, -32'd7207, 32'd414},
{32'd5111, 32'd5918, -32'd7368, 32'd2201},
{32'd12887, 32'd1113, 32'd2744, -32'd21559},
{32'd8674, 32'd664, 32'd103, -32'd12845},
{-32'd7119, -32'd1284, 32'd14114, -32'd4315},
{-32'd8255, 32'd8236, -32'd6115, -32'd11376},
{32'd1445, -32'd2416, -32'd15550, -32'd548},
{32'd10485, 32'd3598, 32'd4354, -32'd8403},
{-32'd7415, -32'd2580, 32'd18064, 32'd1134},
{-32'd2325, -32'd2856, 32'd547, 32'd5259},
{32'd2704, -32'd6667, -32'd5866, -32'd7367},
{-32'd8392, 32'd252, -32'd571, 32'd3204},
{32'd2580, -32'd1323, 32'd4630, -32'd877},
{32'd7949, -32'd486, 32'd4058, -32'd6446},
{-32'd5337, 32'd446, -32'd587, 32'd2222},
{-32'd11921, 32'd12367, 32'd4629, -32'd5713},
{32'd5484, 32'd8667, -32'd3525, -32'd8112},
{32'd406, 32'd109, -32'd8111, 32'd11775},
{32'd2365, 32'd5506, 32'd2757, -32'd11209},
{-32'd2681, 32'd4725, -32'd5613, -32'd1515},
{-32'd3032, -32'd14748, 32'd2563, -32'd1820},
{32'd3274, -32'd5237, 32'd11654, -32'd13587},
{32'd838, -32'd3489, -32'd6510, -32'd7777},
{-32'd186, 32'd12045, 32'd1382, -32'd2360},
{-32'd1621, 32'd12655, 32'd3683, -32'd11339},
{-32'd5857, -32'd6883, -32'd14102, -32'd2953},
{-32'd291, -32'd3834, 32'd5895, -32'd4313},
{-32'd8884, 32'd6517, 32'd6218, 32'd6077},
{-32'd2967, 32'd7719, -32'd3702, 32'd7346},
{-32'd5171, -32'd441, -32'd7425, -32'd5565},
{-32'd1371, 32'd4801, -32'd9989, 32'd7098},
{32'd1276, 32'd11114, 32'd2779, -32'd25000},
{-32'd164, 32'd6085, -32'd3448, -32'd1636},
{-32'd4269, -32'd675, -32'd1225, -32'd13994},
{32'd8777, 32'd12591, 32'd7540, -32'd3074},
{32'd1481, 32'd3754, -32'd8819, 32'd14974},
{-32'd4622, -32'd4150, 32'd10040, -32'd638},
{32'd7966, 32'd14101, -32'd3011, 32'd2812},
{-32'd906, -32'd2207, -32'd7549, -32'd6049},
{32'd14672, -32'd11484, -32'd13391, 32'd1806},
{32'd3326, 32'd4788, 32'd2107, -32'd1132},
{32'd6724, 32'd13537, -32'd936, 32'd2004},
{32'd254, -32'd3594, -32'd6409, -32'd12496},
{32'd11033, 32'd2897, 32'd561, -32'd2595},
{-32'd9522, -32'd660, 32'd11423, 32'd6493},
{-32'd2900, 32'd3042, 32'd12939, -32'd8973},
{32'd6093, 32'd12825, -32'd12381, -32'd3881},
{32'd37, -32'd4485, 32'd4056, 32'd6765},
{-32'd6945, -32'd5810, -32'd3763, -32'd8430},
{-32'd6548, 32'd1349, -32'd3440, -32'd5283},
{32'd1616, 32'd8273, 32'd1720, -32'd3842},
{32'd2240, -32'd4798, -32'd7882, -32'd9886},
{32'd9448, -32'd8541, -32'd20886, -32'd5734},
{-32'd13149, -32'd16042, 32'd12235, -32'd2455},
{32'd9016, -32'd14409, -32'd1995, -32'd3002},
{32'd2721, -32'd4957, 32'd4210, -32'd4228},
{32'd12089, 32'd2047, 32'd11599, 32'd19555},
{32'd4007, 32'd9763, 32'd1019, 32'd6398},
{-32'd7948, 32'd14339, -32'd9692, -32'd4284},
{-32'd748, -32'd807, 32'd561, -32'd5414},
{-32'd6175, -32'd8409, 32'd8294, 32'd3773},
{-32'd6584, 32'd9085, 32'd24540, 32'd27},
{-32'd2289, 32'd8886, 32'd30, 32'd9302},
{-32'd2390, 32'd14466, 32'd9076, 32'd7920},
{-32'd10644, 32'd2559, -32'd9009, 32'd5119},
{-32'd6073, 32'd5232, 32'd12817, -32'd8970},
{-32'd8328, 32'd4123, -32'd13476, 32'd4681},
{-32'd8490, -32'd13715, 32'd6854, -32'd1279},
{-32'd8722, -32'd3643, -32'd1662, 32'd10028},
{-32'd6822, 32'd3916, 32'd3118, 32'd11415},
{-32'd3308, -32'd5100, 32'd5216, -32'd6648},
{-32'd12517, 32'd1575, 32'd670, 32'd8663},
{-32'd12859, 32'd15327, -32'd6721, 32'd7557},
{32'd10156, -32'd14565, -32'd10318, 32'd9209},
{32'd2121, -32'd2369, -32'd351, 32'd14903},
{-32'd10875, -32'd3138, -32'd11283, 32'd9963},
{-32'd1392, 32'd12236, -32'd16272, 32'd2960},
{-32'd3135, -32'd11155, -32'd6891, -32'd3319},
{-32'd15216, 32'd583, 32'd1221, 32'd11145},
{-32'd6334, -32'd2845, -32'd1405, -32'd4149},
{32'd1787, -32'd12278, 32'd7559, -32'd16701},
{-32'd13588, -32'd3362, 32'd230, -32'd1025},
{-32'd135, -32'd1201, 32'd1155, -32'd8755},
{-32'd9058, -32'd2178, 32'd8885, -32'd4965},
{-32'd9704, -32'd62, 32'd4230, -32'd3034},
{-32'd1452, -32'd9690, -32'd488, 32'd3975},
{32'd4113, 32'd979, 32'd11100, 32'd5286},
{-32'd2489, -32'd3317, -32'd17116, 32'd2923},
{-32'd3017, -32'd2436, -32'd7552, 32'd3100},
{32'd4726, 32'd801, 32'd298, 32'd9362},
{32'd8621, -32'd3537, -32'd2589, -32'd14361},
{32'd7519, 32'd4540, -32'd8870, 32'd1904},
{32'd1472, 32'd3801, 32'd676, 32'd8009},
{-32'd2793, 32'd12928, 32'd7907, -32'd12440},
{-32'd10788, -32'd4902, -32'd7546, -32'd4306},
{32'd12817, -32'd63, 32'd4729, -32'd12928},
{-32'd2815, 32'd10315, 32'd12856, -32'd8826},
{32'd8276, 32'd4643, -32'd6598, 32'd8326},
{-32'd4242, 32'd13217, 32'd710, 32'd11399},
{32'd9569, 32'd1192, -32'd15167, -32'd6352},
{-32'd10794, 32'd6515, 32'd7431, -32'd5403},
{-32'd2936, 32'd3325, 32'd12024, -32'd14653},
{-32'd950, -32'd9545, 32'd5216, 32'd9538},
{-32'd7354, 32'd321, 32'd8607, -32'd4118},
{32'd12203, 32'd6337, -32'd7190, -32'd954},
{-32'd5824, -32'd10743, 32'd2405, -32'd5991},
{32'd8726, 32'd5218, 32'd12590, -32'd2874},
{-32'd2353, -32'd9624, 32'd2199, 32'd3062},
{-32'd6031, 32'd4154, 32'd2496, -32'd1181},
{-32'd16065, -32'd2720, -32'd5631, 32'd9341},
{32'd11156, 32'd4284, 32'd2931, 32'd7043},
{-32'd10038, 32'd12191, 32'd2915, 32'd5164},
{32'd10002, 32'd10399, 32'd12108, 32'd10659},
{32'd4226, 32'd9638, -32'd3075, 32'd4988},
{32'd3513, 32'd5183, 32'd1634, 32'd10626},
{32'd1221, 32'd3435, 32'd7810, 32'd6876},
{-32'd310, 32'd2939, -32'd14137, -32'd2534},
{-32'd11547, 32'd1072, -32'd4770, 32'd3364},
{-32'd9743, -32'd15838, 32'd255, -32'd616},
{-32'd11197, 32'd1996, 32'd8909, 32'd384},
{-32'd3580, -32'd11699, -32'd5717, 32'd4066},
{32'd6684, -32'd4811, -32'd7403, 32'd7816},
{32'd5224, 32'd8874, -32'd2012, -32'd2133},
{32'd1276, 32'd1040, 32'd7510, 32'd3772},
{32'd10122, 32'd4497, -32'd2728, 32'd10031},
{-32'd4914, 32'd2692, -32'd3580, 32'd6554},
{-32'd5761, 32'd12473, -32'd250, 32'd3409},
{32'd2175, -32'd7787, 32'd5445, 32'd10880},
{32'd905, 32'd2341, -32'd6641, -32'd313},
{-32'd3994, -32'd6534, -32'd7639, 32'd5583},
{32'd6857, 32'd11928, 32'd3172, -32'd10201},
{-32'd5151, 32'd4320, -32'd12355, 32'd898},
{-32'd1187, 32'd1696, -32'd783, 32'd9059},
{32'd3427, 32'd7816, -32'd1030, -32'd2373},
{32'd9917, -32'd10973, 32'd3078, 32'd1690},
{-32'd4324, -32'd16400, -32'd1566, 32'd4812},
{32'd173, -32'd3781, -32'd1585, 32'd2862},
{-32'd2235, 32'd7233, -32'd10258, 32'd1145},
{-32'd3853, -32'd844, 32'd1389, 32'd1102},
{32'd4016, 32'd515, -32'd9591, 32'd6623},
{-32'd6943, 32'd6253, 32'd1041, -32'd8204},
{-32'd5688, 32'd4135, 32'd12254, -32'd10099},
{-32'd401, 32'd803, 32'd10677, -32'd6723},
{32'd7025, -32'd1191, 32'd11951, 32'd5469},
{32'd8405, -32'd3499, 32'd7648, -32'd5644},
{-32'd7968, -32'd785, 32'd11450, -32'd16225},
{32'd11643, 32'd5115, -32'd9050, -32'd7171},
{32'd4352, 32'd6219, -32'd10681, 32'd1746},
{32'd3385, -32'd9221, -32'd4577, -32'd9946},
{-32'd6915, -32'd866, 32'd1837, -32'd7953},
{32'd6370, -32'd768, 32'd2393, 32'd6689},
{-32'd272, -32'd4508, 32'd8777, 32'd134},
{32'd5909, 32'd3317, -32'd5612, -32'd7058},
{-32'd2390, 32'd5984, -32'd3150, -32'd8953},
{32'd13178, 32'd2275, 32'd3004, 32'd4322},
{-32'd6821, 32'd1234, 32'd922, -32'd12403},
{32'd2686, 32'd3475, 32'd10643, 32'd12821},
{32'd2233, 32'd655, 32'd420, -32'd6501},
{32'd3805, 32'd2590, 32'd6462, -32'd672},
{32'd2767, -32'd1013, -32'd6609, -32'd8807},
{-32'd2671, 32'd6380, -32'd12970, 32'd5338},
{32'd3935, -32'd10701, -32'd4213, -32'd10848},
{32'd9996, -32'd11254, -32'd12033, -32'd6556},
{32'd4958, -32'd9386, 32'd5720, -32'd12280},
{-32'd3476, 32'd7561, 32'd4681, 32'd1124},
{-32'd8643, -32'd4137, -32'd9409, -32'd1088},
{32'd5346, -32'd4802, 32'd4545, -32'd12798},
{-32'd12114, -32'd3897, 32'd2050, 32'd453},
{32'd6320, -32'd11201, -32'd14890, 32'd8742},
{-32'd5956, -32'd4746, -32'd5844, 32'd5757},
{32'd6176, 32'd2077, -32'd2869, 32'd5763},
{32'd12879, 32'd9211, -32'd13875, 32'd7002},
{-32'd10364, 32'd3004, -32'd3430, 32'd11714},
{-32'd9205, -32'd4585, 32'd4261, 32'd11143},
{-32'd6803, -32'd9607, 32'd6865, -32'd3755},
{-32'd8941, 32'd1427, 32'd13081, 32'd3362},
{32'd10754, -32'd12252, 32'd3393, 32'd7300},
{-32'd2158, -32'd406, 32'd10654, 32'd3835},
{32'd1111, 32'd3021, 32'd1727, 32'd7104},
{32'd3412, 32'd3554, 32'd6713, -32'd5009},
{-32'd6198, 32'd1289, 32'd3562, -32'd5252},
{32'd5587, 32'd3527, 32'd6170, -32'd5788},
{32'd6532, 32'd3631, 32'd1212, 32'd5419},
{-32'd546, -32'd7578, -32'd3246, 32'd5509},
{-32'd11654, -32'd291, -32'd9031, -32'd3470},
{32'd1548, 32'd14910, -32'd4467, 32'd6772},
{32'd10378, -32'd1419, 32'd613, -32'd1304},
{-32'd5874, 32'd2225, 32'd14877, -32'd4013},
{32'd453, -32'd4176, 32'd6415, 32'd2157},
{-32'd5393, 32'd3784, -32'd2203, 32'd16962},
{-32'd367, -32'd3492, 32'd3810, 32'd7794},
{-32'd8339, 32'd2129, -32'd297, -32'd18227},
{-32'd8958, 32'd3754, 32'd16704, -32'd10356},
{32'd8135, 32'd4208, 32'd17700, -32'd9600},
{-32'd4672, 32'd7791, 32'd12771, -32'd4389},
{-32'd4385, -32'd2192, -32'd3301, 32'd4092},
{-32'd10444, -32'd4991, -32'd7605, -32'd5025},
{-32'd2113, 32'd1707, 32'd9365, 32'd11420},
{-32'd4301, -32'd3554, -32'd4775, 32'd5593},
{-32'd1137, -32'd11523, -32'd5999, -32'd4360},
{-32'd3230, -32'd10925, 32'd8185, -32'd1698},
{-32'd2376, 32'd576, -32'd2829, 32'd2706},
{32'd3523, -32'd3641, 32'd650, -32'd11811},
{32'd1526, -32'd5048, 32'd2694, -32'd5537},
{32'd1504, -32'd1598, -32'd6834, 32'd7972},
{-32'd4330, -32'd4640, 32'd348, -32'd7071},
{-32'd7263, 32'd1168, -32'd8574, -32'd171},
{-32'd2661, 32'd1726, 32'd11522, -32'd13874},
{32'd4005, -32'd12071, -32'd9833, -32'd4614},
{-32'd10867, -32'd4054, 32'd7992, 32'd1325},
{-32'd3097, 32'd3861, 32'd15140, -32'd8921},
{-32'd4193, -32'd5976, 32'd1203, 32'd7064},
{-32'd15747, 32'd3929, 32'd7982, 32'd2163},
{-32'd8899, -32'd2185, -32'd2648, -32'd11474},
{32'd10417, 32'd6167, -32'd502, 32'd3807},
{-32'd2593, 32'd6043, 32'd2833, -32'd420},
{-32'd113, -32'd4674, -32'd2107, 32'd144},
{32'd1865, -32'd1167, 32'd9397, 32'd12379},
{32'd10534, 32'd10101, -32'd9839, 32'd2115},
{-32'd3423, -32'd3499, 32'd3270, 32'd704},
{-32'd2535, -32'd7165, 32'd16443, 32'd14212},
{-32'd10336, 32'd109, 32'd99, 32'd4783},
{-32'd3566, 32'd4814, 32'd10886, -32'd7760},
{-32'd18398, -32'd2933, 32'd8059, -32'd3680},
{32'd1973, -32'd2272, -32'd2961, 32'd853},
{-32'd5433, 32'd14493, 32'd6643, -32'd13161},
{32'd4742, 32'd2060, -32'd4920, -32'd1182},
{-32'd231, -32'd7518, -32'd13586, -32'd1748},
{32'd8341, 32'd456, -32'd9886, 32'd4459},
{32'd5808, 32'd1394, -32'd8068, 32'd12568},
{32'd3444, -32'd458, -32'd3213, -32'd12121},
{-32'd2095, 32'd2246, -32'd14010, 32'd7176},
{32'd794, -32'd9818, 32'd1244, 32'd6305},
{32'd2500, 32'd1074, -32'd2938, -32'd2271},
{32'd4131, 32'd9081, -32'd2409, -32'd5974},
{32'd13459, 32'd2440, -32'd2624, -32'd5374},
{32'd6350, -32'd893, 32'd12688, 32'd10315},
{-32'd20498, -32'd8799, -32'd10117, 32'd1012}
},
{{32'd5628, 32'd16548, 32'd8750, 32'd1887},
{-32'd12599, -32'd8069, 32'd1655, 32'd959},
{-32'd2649, -32'd7345, 32'd18079, -32'd3839},
{32'd4503, 32'd12380, 32'd195, 32'd1872},
{32'd2160, -32'd10052, -32'd5138, -32'd3058},
{-32'd5571, -32'd6448, -32'd17249, -32'd12719},
{32'd2067, -32'd1444, -32'd257, -32'd8463},
{32'd10350, -32'd3315, -32'd2057, -32'd13260},
{-32'd5527, 32'd2570, 32'd885, 32'd4380},
{32'd16714, 32'd11757, 32'd3315, -32'd1493},
{-32'd13139, -32'd4780, 32'd5379, -32'd4759},
{-32'd5525, -32'd6053, -32'd6217, -32'd8439},
{-32'd8652, 32'd7068, 32'd4146, -32'd2202},
{-32'd6045, 32'd1301, 32'd6037, -32'd6227},
{-32'd3942, 32'd4600, 32'd3225, 32'd2112},
{-32'd11147, -32'd3592, 32'd11191, -32'd4818},
{32'd6446, 32'd7610, 32'd441, 32'd4753},
{-32'd8769, 32'd4120, 32'd19329, 32'd11353},
{32'd1325, 32'd669, -32'd2784, -32'd1144},
{-32'd0, -32'd1788, 32'd69, 32'd377},
{-32'd3854, 32'd2441, 32'd5826, -32'd2155},
{-32'd3750, -32'd1976, 32'd2392, -32'd9430},
{-32'd4810, -32'd380, 32'd3076, -32'd4767},
{32'd3457, -32'd8318, 32'd1991, 32'd3035},
{32'd9832, 32'd3793, -32'd2629, -32'd5941},
{32'd10909, 32'd5320, -32'd10827, -32'd5386},
{32'd5842, 32'd5900, -32'd1206, 32'd1265},
{32'd12, 32'd3538, -32'd2739, -32'd752},
{32'd957, 32'd7961, 32'd5063, 32'd2916},
{-32'd401, 32'd3041, -32'd4036, 32'd2693},
{32'd8701, -32'd623, -32'd16191, -32'd7160},
{32'd2744, -32'd4136, -32'd1423, 32'd969},
{32'd4283, -32'd636, -32'd2375, 32'd875},
{-32'd8849, -32'd9136, -32'd5004, -32'd7411},
{32'd10564, 32'd8200, 32'd557, 32'd4190},
{-32'd8536, -32'd3887, 32'd17005, 32'd7270},
{32'd2964, -32'd3410, -32'd8383, -32'd3356},
{-32'd2259, -32'd5263, 32'd740, 32'd4654},
{-32'd8942, 32'd637, 32'd1146, -32'd1377},
{-32'd1840, -32'd4302, -32'd3109, -32'd1899},
{32'd4532, 32'd790, -32'd7494, -32'd4586},
{32'd8887, 32'd11441, 32'd13827, -32'd2669},
{-32'd2355, 32'd5019, 32'd10670, 32'd5063},
{-32'd10178, -32'd9875, -32'd10873, -32'd4039},
{32'd7196, -32'd3743, -32'd5824, 32'd7090},
{-32'd1434, -32'd442, -32'd11770, -32'd2105},
{32'd6366, -32'd4279, 32'd4092, 32'd4062},
{-32'd4214, -32'd14655, -32'd13153, 32'd5060},
{-32'd5652, 32'd8639, 32'd11543, -32'd561},
{32'd7312, 32'd1689, -32'd2345, 32'd1902},
{32'd1417, -32'd5486, -32'd7655, 32'd7377},
{32'd3705, 32'd6672, 32'd5948, 32'd210},
{32'd1989, -32'd1792, 32'd6311, -32'd1142},
{-32'd1649, -32'd2148, 32'd5835, 32'd9541},
{32'd14092, -32'd699, 32'd3877, -32'd1569},
{-32'd1836, 32'd567, -32'd11380, -32'd8314},
{-32'd10597, 32'd433, -32'd1916, 32'd3406},
{-32'd885, -32'd1358, 32'd3998, 32'd12710},
{32'd1116, -32'd2434, 32'd384, -32'd6609},
{-32'd1705, -32'd3475, -32'd7848, -32'd3815},
{-32'd8146, -32'd13090, -32'd10350, -32'd6144},
{-32'd797, 32'd2035, 32'd1448, -32'd9230},
{-32'd7835, -32'd5490, -32'd44, 32'd3296},
{-32'd4980, 32'd5544, -32'd887, -32'd6460},
{-32'd7560, -32'd2289, -32'd222, 32'd2624},
{32'd5505, 32'd6162, 32'd8871, 32'd7692},
{32'd3805, 32'd4189, -32'd12538, -32'd8031},
{-32'd5335, -32'd5119, -32'd2500, 32'd857},
{-32'd2746, -32'd2737, 32'd4850, 32'd391},
{32'd11280, -32'd6598, -32'd2652, 32'd348},
{32'd1565, -32'd5290, -32'd4794, -32'd4512},
{-32'd3887, -32'd7884, 32'd3678, -32'd6672},
{-32'd1999, -32'd3384, -32'd2909, -32'd533},
{-32'd1562, -32'd1335, -32'd6586, -32'd6190},
{32'd3022, 32'd1527, -32'd4305, -32'd401},
{-32'd7019, -32'd8219, 32'd7867, 32'd7369},
{32'd3366, -32'd4900, -32'd5557, 32'd7329},
{-32'd3684, 32'd2422, -32'd347, -32'd3311},
{-32'd6483, 32'd1826, 32'd1189, 32'd16738},
{-32'd1637, 32'd1409, 32'd5643, 32'd10675},
{32'd18598, 32'd9537, 32'd2696, 32'd637},
{32'd5733, 32'd3228, 32'd10360, 32'd4830},
{-32'd16327, -32'd6741, -32'd4851, -32'd5781},
{-32'd8555, 32'd53, -32'd2649, 32'd2906},
{-32'd11571, -32'd2089, 32'd5, 32'd5304},
{32'd1896, 32'd6929, 32'd613, -32'd8379},
{-32'd2045, -32'd6071, 32'd4330, 32'd2570},
{-32'd11196, -32'd7220, 32'd879, -32'd8380},
{-32'd11361, -32'd2473, -32'd5609, 32'd427},
{32'd469, -32'd5221, 32'd3608, -32'd3507},
{32'd10334, 32'd1182, -32'd1247, -32'd7643},
{-32'd10533, -32'd2452, 32'd6026, 32'd2873},
{32'd4863, 32'd8956, 32'd12644, -32'd498},
{32'd911, 32'd3606, 32'd2483, 32'd2301},
{32'd8805, -32'd1311, 32'd9935, 32'd9482},
{32'd8859, 32'd4795, -32'd11379, 32'd3247},
{32'd12464, 32'd6362, 32'd1017, -32'd1881},
{32'd6814, -32'd1034, 32'd9272, 32'd3112},
{-32'd4636, -32'd2157, 32'd613, 32'd5382},
{32'd6429, 32'd11983, 32'd5882, 32'd2575},
{32'd411, 32'd772, 32'd812, 32'd796},
{32'd7013, 32'd1777, 32'd7417, -32'd7023},
{32'd226, -32'd8980, -32'd4833, -32'd2665},
{-32'd5422, 32'd3105, -32'd2087, 32'd1462},
{-32'd4591, 32'd3503, 32'd472, 32'd7351},
{32'd7805, -32'd3572, 32'd1072, -32'd2530},
{-32'd13488, -32'd73, -32'd2450, 32'd3341},
{32'd3997, -32'd6674, -32'd2187, -32'd18962},
{32'd9323, 32'd4756, 32'd773, 32'd5935},
{32'd3907, 32'd1075, -32'd8578, 32'd4146},
{-32'd9089, -32'd7959, 32'd6175, 32'd5753},
{32'd2295, 32'd3697, 32'd7476, -32'd1556},
{-32'd1172, 32'd2349, 32'd4361, 32'd1022},
{32'd350, 32'd669, 32'd3707, -32'd6852},
{-32'd2201, -32'd3032, -32'd8424, 32'd1802},
{-32'd11782, -32'd3986, -32'd5812, -32'd2789},
{-32'd8422, 32'd1086, -32'd3234, -32'd4604},
{32'd10472, -32'd3203, 32'd316, 32'd5843},
{32'd440, -32'd7886, -32'd2678, -32'd815},
{32'd12260, 32'd10063, 32'd5491, 32'd5077},
{-32'd7534, 32'd9191, 32'd15553, -32'd4489},
{-32'd4595, 32'd3449, 32'd10423, 32'd108},
{-32'd1412, 32'd1704, -32'd793, -32'd11311},
{32'd9622, -32'd1652, 32'd4113, 32'd2976},
{-32'd2743, 32'd1755, 32'd5722, 32'd5288},
{32'd12737, -32'd793, -32'd604, -32'd9464},
{-32'd7090, 32'd966, 32'd3337, -32'd2522},
{32'd636, -32'd3887, 32'd1737, 32'd2978},
{-32'd511, -32'd11899, -32'd7911, -32'd13710},
{-32'd3522, -32'd1503, -32'd2337, -32'd11019},
{-32'd7703, -32'd2486, 32'd13309, -32'd1811},
{32'd7495, -32'd11716, -32'd8338, -32'd2506},
{-32'd3273, -32'd12594, -32'd12563, -32'd1954},
{32'd4022, 32'd2007, -32'd2511, -32'd6452},
{32'd3035, 32'd9822, 32'd2859, 32'd3807},
{32'd912, 32'd9772, 32'd9529, -32'd5542},
{-32'd1661, 32'd4381, 32'd1120, 32'd12912},
{32'd6220, 32'd3253, -32'd1485, 32'd2948},
{-32'd4330, 32'd7557, 32'd12671, -32'd5325},
{32'd2837, -32'd6023, -32'd4148, 32'd518},
{32'd10871, 32'd420, -32'd4880, 32'd5272},
{32'd1192, 32'd1137, 32'd1549, -32'd1661},
{-32'd528, 32'd5097, 32'd7768, -32'd2361},
{32'd242, 32'd4645, -32'd3345, -32'd2805},
{-32'd7960, 32'd4939, 32'd1717, -32'd2431},
{32'd3523, 32'd2543, 32'd4376, 32'd346},
{-32'd13098, -32'd3946, 32'd889, -32'd2022},
{-32'd6928, -32'd4397, 32'd3355, 32'd0},
{32'd158, -32'd2067, -32'd268, -32'd1619},
{-32'd444, -32'd3683, -32'd4068, -32'd5270},
{-32'd12009, -32'd2502, -32'd623, -32'd160},
{32'd12418, 32'd7792, -32'd2280, 32'd5985},
{-32'd5824, 32'd2541, 32'd5516, 32'd6501},
{32'd4959, -32'd1498, -32'd5605, -32'd3727},
{-32'd8658, -32'd10204, -32'd9302, -32'd336},
{32'd6152, 32'd4173, 32'd6143, 32'd10303},
{32'd1840, 32'd7096, -32'd822, 32'd9569},
{32'd2980, 32'd4082, -32'd1867, 32'd3117},
{-32'd8925, 32'd7863, 32'd9608, -32'd122},
{32'd2758, 32'd1131, 32'd4921, 32'd602},
{-32'd7819, 32'd731, 32'd5452, 32'd1490},
{32'd4204, 32'd5724, 32'd4922, 32'd1331},
{-32'd15645, -32'd5353, 32'd6528, -32'd15744},
{32'd4491, 32'd196, 32'd6014, -32'd2597},
{32'd5384, 32'd446, 32'd2627, 32'd11333},
{32'd1796, -32'd11040, -32'd7526, -32'd697},
{32'd8274, -32'd307, -32'd1002, 32'd14634},
{-32'd10886, -32'd7943, 32'd190, 32'd4491},
{-32'd4429, -32'd7648, -32'd935, 32'd5204},
{-32'd13083, -32'd10483, -32'd2096, 32'd680},
{-32'd2074, -32'd10997, -32'd5068, -32'd3699},
{32'd1029, -32'd2707, -32'd13010, -32'd1580},
{32'd12454, 32'd4835, -32'd3215, -32'd1640},
{-32'd5355, -32'd1131, 32'd28, -32'd2592},
{32'd4927, 32'd2523, -32'd6976, -32'd2515},
{32'd1058, -32'd3618, -32'd9181, -32'd4260},
{32'd15212, -32'd6223, -32'd14539, 32'd2934},
{-32'd9377, 32'd1179, -32'd3085, -32'd3436},
{32'd3076, 32'd4007, 32'd7286, 32'd415},
{-32'd13441, -32'd3146, -32'd7960, -32'd5021},
{-32'd1824, -32'd5250, 32'd7029, 32'd1819},
{-32'd7277, 32'd898, -32'd625, -32'd1991},
{32'd2931, 32'd935, -32'd3991, -32'd4739},
{32'd120, -32'd5443, -32'd463, -32'd7221},
{-32'd7889, -32'd601, -32'd2915, 32'd7075},
{32'd3184, 32'd4159, -32'd6681, -32'd11131},
{32'd4980, 32'd8584, 32'd5464, 32'd5344},
{-32'd13134, -32'd3804, 32'd6361, -32'd1650},
{-32'd13011, -32'd2910, -32'd5518, 32'd1284},
{-32'd5651, 32'd850, 32'd3836, -32'd1262},
{-32'd3562, 32'd2450, 32'd3943, 32'd1343},
{32'd2661, -32'd10119, -32'd283, 32'd7858},
{-32'd612, -32'd1226, -32'd6459, 32'd6718},
{32'd12647, 32'd8688, 32'd4648, -32'd1189},
{-32'd716, -32'd5860, 32'd5346, -32'd8467},
{32'd6947, 32'd10903, 32'd3754, -32'd8001},
{-32'd2311, -32'd1389, -32'd9943, 32'd1954},
{32'd1065, 32'd2422, 32'd1058, -32'd12160},
{-32'd4900, -32'd3609, -32'd8980, -32'd612},
{32'd11477, 32'd5057, 32'd3663, 32'd1651},
{-32'd9175, -32'd5379, -32'd5576, 32'd1760},
{32'd5163, 32'd2728, -32'd435, -32'd11619},
{-32'd9661, -32'd7888, -32'd7167, -32'd1447},
{32'd164, -32'd842, -32'd11522, 32'd10567},
{-32'd7591, -32'd8987, -32'd2833, 32'd146},
{32'd7704, 32'd3548, -32'd6425, 32'd9524},
{-32'd5707, -32'd659, -32'd3, -32'd5294},
{32'd4855, -32'd4170, -32'd9561, -32'd2434},
{32'd9133, -32'd4744, 32'd2842, 32'd8831},
{32'd504, 32'd1193, 32'd8544, 32'd2554},
{-32'd10842, -32'd6187, -32'd10500, 32'd1841},
{-32'd16429, 32'd379, 32'd1130, -32'd3057},
{-32'd8030, -32'd1228, 32'd11073, 32'd3243},
{32'd5465, -32'd984, 32'd3945, 32'd5213},
{32'd9225, 32'd928, -32'd6992, -32'd5691},
{-32'd14009, 32'd1604, 32'd909, 32'd5824},
{32'd4028, -32'd9321, -32'd10666, -32'd1893},
{-32'd3229, -32'd4797, -32'd12362, 32'd5196},
{32'd5331, -32'd2263, -32'd2583, -32'd13033},
{-32'd1168, -32'd1394, 32'd8818, 32'd13330},
{-32'd6294, -32'd6056, 32'd3605, 32'd2395},
{-32'd2828, 32'd1652, 32'd9323, 32'd8630},
{32'd2892, 32'd6448, 32'd11710, -32'd3148},
{-32'd5196, -32'd1268, 32'd3728, -32'd7462},
{-32'd10686, 32'd2297, 32'd1526, -32'd7792},
{-32'd11357, -32'd8464, -32'd920, 32'd3006},
{32'd6470, -32'd2552, -32'd3066, 32'd3942},
{-32'd3776, 32'd1396, 32'd1743, -32'd12598},
{32'd7261, 32'd7789, 32'd14014, 32'd6375},
{-32'd633, -32'd1062, -32'd1921, 32'd6002},
{-32'd3342, -32'd3200, 32'd4756, 32'd9540},
{-32'd6782, -32'd4792, -32'd5745, 32'd636},
{-32'd6129, 32'd6180, 32'd5652, -32'd9425},
{32'd7768, 32'd4182, 32'd6584, -32'd425},
{32'd879, -32'd4178, -32'd4449, 32'd186},
{-32'd6929, -32'd2672, -32'd764, 32'd228},
{-32'd5876, -32'd10815, -32'd116, -32'd390},
{32'd325, 32'd2172, -32'd9469, -32'd1640},
{32'd6824, 32'd8877, 32'd2375, -32'd1099},
{-32'd6351, -32'd5550, 32'd5704, -32'd180},
{-32'd9867, 32'd6589, 32'd13824, 32'd3485},
{32'd658, -32'd1686, 32'd4344, 32'd6516},
{-32'd6155, -32'd7844, -32'd6519, -32'd8226},
{-32'd4730, 32'd482, -32'd5033, 32'd10311},
{32'd11474, 32'd13472, 32'd2486, 32'd3719},
{32'd10002, -32'd374, -32'd11741, -32'd821},
{32'd4903, -32'd8857, -32'd725, 32'd5804},
{-32'd1185, 32'd6315, -32'd3561, -32'd3527},
{-32'd1032, -32'd6079, 32'd3954, 32'd24},
{-32'd11454, -32'd754, -32'd5868, -32'd2716},
{32'd1202, -32'd1396, 32'd1723, 32'd8547},
{32'd2999, -32'd185, -32'd5390, 32'd6982},
{32'd7466, 32'd2310, -32'd8717, 32'd1010},
{-32'd5325, -32'd877, 32'd3891, -32'd8910},
{32'd1944, -32'd7576, 32'd2044, -32'd5848},
{32'd7898, -32'd4281, 32'd9288, 32'd7208},
{32'd11366, 32'd911, -32'd6406, -32'd7857},
{32'd7480, 32'd1738, -32'd6212, 32'd486},
{-32'd7429, -32'd2490, -32'd1959, 32'd3055},
{32'd2859, -32'd6868, -32'd520, -32'd9764},
{-32'd8157, -32'd178, -32'd4751, -32'd1405},
{-32'd16082, -32'd856, 32'd1874, 32'd335},
{-32'd546, -32'd7655, 32'd6910, 32'd8663},
{32'd4043, -32'd4722, 32'd5521, 32'd5329},
{-32'd4058, 32'd223, -32'd5650, 32'd11112},
{32'd8573, 32'd2584, 32'd13924, -32'd3866},
{-32'd6701, 32'd1034, -32'd1030, 32'd12410},
{32'd2807, 32'd127, 32'd13627, 32'd4409},
{-32'd9347, -32'd6818, 32'd3707, 32'd1194},
{-32'd5371, -32'd6746, 32'd9120, 32'd8347},
{32'd8920, 32'd4273, -32'd9662, 32'd5058},
{-32'd8030, -32'd2199, -32'd2323, 32'd10130},
{-32'd1429, -32'd4752, 32'd1848, 32'd9079},
{-32'd11851, -32'd8650, -32'd4227, -32'd8673},
{-32'd2094, -32'd8579, 32'd5273, 32'd3147},
{-32'd16425, 32'd94, -32'd1342, -32'd9887},
{32'd13595, 32'd12700, 32'd5676, 32'd1965},
{-32'd2935, 32'd4517, -32'd3574, 32'd2357},
{-32'd8477, -32'd5587, -32'd7522, -32'd5124},
{-32'd183, -32'd989, -32'd5060, -32'd8490},
{32'd3741, 32'd7666, 32'd3546, -32'd3938},
{-32'd6916, -32'd27, -32'd175, 32'd3136},
{32'd138, 32'd7525, -32'd2327, 32'd418},
{-32'd4673, -32'd865, -32'd5438, -32'd3484},
{32'd12441, -32'd160, 32'd2716, -32'd4770},
{32'd8358, -32'd15002, -32'd3293, 32'd1205},
{32'd1861, -32'd1862, -32'd2986, 32'd2223},
{32'd6421, -32'd876, 32'd906, 32'd7495},
{-32'd17094, -32'd2454, -32'd1800, -32'd5090},
{32'd8691, 32'd4884, 32'd10927, -32'd4915},
{32'd5514, 32'd7722, 32'd5973, -32'd1209},
{-32'd2692, 32'd3381, 32'd1045, -32'd2211},
{32'd23501, 32'd8822, -32'd7306, 32'd5640},
{-32'd1994, 32'd4218, 32'd6062, -32'd273},
{32'd4754, -32'd3914, -32'd4853, -32'd860},
{32'd6163, -32'd6319, -32'd3559, -32'd4632},
{-32'd12313, -32'd2411, 32'd9195, 32'd7489},
{-32'd3294, 32'd11566, 32'd8963, 32'd7652},
{32'd5464, 32'd4825, -32'd7973, -32'd8491},
{-32'd8755, -32'd1747, 32'd6310, -32'd5068}
},
{{32'd5678, 32'd12463, -32'd4524, 32'd7028},
{-32'd4108, -32'd9579, 32'd6699, -32'd3221},
{32'd8075, -32'd1661, 32'd2424, 32'd3920},
{32'd3909, -32'd6389, 32'd569, 32'd2402},
{-32'd13209, 32'd3896, -32'd6903, 32'd2405},
{32'd4687, 32'd1767, -32'd5781, 32'd5985},
{-32'd1013, 32'd8643, 32'd5556, 32'd12613},
{32'd650, -32'd217, 32'd5395, 32'd12551},
{-32'd7844, 32'd6032, 32'd5337, -32'd5382},
{32'd8678, 32'd8798, 32'd4836, 32'd9433},
{32'd2877, 32'd2556, -32'd2154, -32'd4132},
{-32'd1067, 32'd2917, 32'd2178, -32'd4030},
{-32'd5912, -32'd4300, 32'd10605, 32'd9638},
{-32'd4105, -32'd105, 32'd1765, 32'd1557},
{-32'd13359, -32'd10398, 32'd7255, -32'd4957},
{32'd4785, -32'd6551, -32'd571, 32'd4015},
{32'd2196, 32'd159, -32'd442, 32'd8116},
{32'd8128, 32'd5126, 32'd6254, -32'd4858},
{-32'd1612, -32'd6329, 32'd4767, -32'd1953},
{32'd2504, 32'd6294, 32'd1761, -32'd3700},
{-32'd4025, -32'd9889, -32'd7572, -32'd6170},
{-32'd1036, -32'd471, -32'd1829, -32'd13368},
{-32'd5844, -32'd11001, -32'd902, 32'd17478},
{32'd861, -32'd13432, -32'd891, -32'd7241},
{32'd4848, 32'd6926, -32'd1248, 32'd7390},
{32'd12676, 32'd2858, 32'd7179, -32'd3216},
{32'd923, -32'd5879, -32'd7389, -32'd4318},
{-32'd5072, 32'd1788, 32'd10560, 32'd17701},
{32'd5024, -32'd9736, 32'd853, -32'd9196},
{-32'd8916, 32'd6841, 32'd9116, 32'd131},
{32'd6675, 32'd3120, 32'd4872, 32'd14392},
{32'd3046, -32'd4515, -32'd9243, -32'd8589},
{32'd4718, 32'd4618, 32'd4418, 32'd14396},
{-32'd9030, -32'd1028, -32'd6356, -32'd5085},
{32'd2839, 32'd9957, 32'd9541, 32'd5109},
{-32'd1284, 32'd3296, -32'd1019, -32'd851},
{-32'd7795, 32'd195, 32'd7916, 32'd2153},
{32'd3461, -32'd112, 32'd2989, 32'd734},
{32'd814, 32'd3314, 32'd8556, 32'd6943},
{-32'd2728, 32'd1584, 32'd16592, -32'd3005},
{-32'd4190, -32'd8985, -32'd3196, -32'd7440},
{32'd13984, 32'd729, 32'd15676, 32'd4734},
{-32'd6853, 32'd4039, 32'd4755, -32'd6442},
{-32'd8393, -32'd2076, 32'd5606, 32'd1473},
{-32'd3291, 32'd1569, -32'd12879, 32'd8398},
{-32'd344, 32'd5330, 32'd14984, -32'd6524},
{32'd2188, 32'd3441, -32'd6213, -32'd4856},
{32'd5891, -32'd7499, -32'd7860, -32'd4303},
{32'd6676, 32'd1368, -32'd5997, 32'd3537},
{32'd391, -32'd6223, 32'd2486, 32'd1137},
{-32'd12431, 32'd2125, 32'd972, 32'd6860},
{-32'd4924, -32'd2973, -32'd8086, -32'd5913},
{32'd629, -32'd5879, 32'd7122, -32'd8583},
{-32'd282, 32'd1970, -32'd6227, -32'd2899},
{-32'd16535, -32'd11588, -32'd2034, -32'd4459},
{32'd4741, -32'd696, 32'd3301, 32'd4704},
{32'd6674, 32'd2223, 32'd4114, 32'd2302},
{-32'd14419, -32'd10341, 32'd341, 32'd5644},
{32'd2119, 32'd1006, 32'd915, -32'd4511},
{32'd3842, -32'd1985, 32'd2720, -32'd3341},
{-32'd3637, 32'd3433, -32'd3219, 32'd1843},
{-32'd9319, 32'd5410, 32'd8960, 32'd2202},
{-32'd6364, -32'd14102, 32'd471, -32'd7095},
{32'd4404, -32'd2859, -32'd1481, -32'd4962},
{-32'd9847, -32'd173, 32'd2716, 32'd12686},
{-32'd6012, 32'd8864, 32'd14618, 32'd8064},
{32'd3167, 32'd1571, 32'd1074, 32'd3186},
{32'd3388, -32'd6725, 32'd9047, 32'd6018},
{-32'd567, -32'd6490, 32'd4162, -32'd8959},
{-32'd6891, 32'd2089, 32'd5502, -32'd8},
{-32'd3047, -32'd5345, -32'd1549, 32'd8767},
{-32'd1879, 32'd3041, -32'd3603, 32'd386},
{32'd448, 32'd2812, -32'd1407, -32'd5611},
{32'd5168, -32'd17349, 32'd7316, -32'd1709},
{-32'd7856, 32'd2855, 32'd3223, 32'd2055},
{-32'd5610, 32'd1895, 32'd6954, -32'd656},
{-32'd6645, -32'd4654, -32'd7596, -32'd1383},
{32'd2139, -32'd1640, 32'd1773, 32'd5676},
{-32'd5118, 32'd13887, 32'd10815, -32'd4175},
{32'd2245, 32'd1702, 32'd289, -32'd5905},
{32'd754, 32'd2812, -32'd6689, -32'd3467},
{32'd6342, 32'd5467, 32'd330, -32'd2020},
{-32'd7261, -32'd2072, -32'd6702, -32'd3776},
{32'd8122, -32'd10439, -32'd16353, -32'd4487},
{-32'd9797, -32'd3633, -32'd9954, 32'd6674},
{32'd8223, -32'd9643, -32'd3244, -32'd4627},
{-32'd11505, -32'd4378, 32'd2252, 32'd189},
{-32'd6340, -32'd14701, 32'd2003, -32'd4412},
{-32'd1805, 32'd2685, -32'd132, -32'd2768},
{-32'd5922, -32'd5067, -32'd4700, -32'd8821},
{32'd4391, 32'd1904, 32'd12775, 32'd2222},
{32'd237, -32'd7913, 32'd9510, 32'd2727},
{-32'd927, 32'd15696, 32'd2112, 32'd10026},
{-32'd4539, -32'd902, 32'd7902, 32'd6798},
{-32'd990, -32'd1075, 32'd8093, -32'd7095},
{-32'd2865, -32'd970, -32'd1149, 32'd1639},
{-32'd3453, 32'd8107, -32'd3382, 32'd6835},
{32'd83, 32'd12104, 32'd45, 32'd13151},
{32'd4334, -32'd1994, 32'd12333, -32'd1398},
{32'd5485, 32'd9427, -32'd1437, 32'd3222},
{-32'd6967, 32'd1880, -32'd7805, -32'd13283},
{-32'd2842, -32'd340, -32'd8471, 32'd9796},
{32'd5936, 32'd15136, -32'd4772, -32'd7793},
{32'd2634, -32'd2393, -32'd4405, 32'd4996},
{32'd2914, 32'd2572, 32'd6986, 32'd5427},
{-32'd5205, 32'd104, -32'd4471, 32'd4514},
{32'd10843, 32'd2998, -32'd2771, -32'd8199},
{32'd4988, -32'd3882, -32'd3818, 32'd2103},
{32'd355, -32'd5129, -32'd9561, -32'd5926},
{-32'd2429, -32'd5320, -32'd5240, 32'd1903},
{-32'd9145, 32'd1058, -32'd6643, 32'd8699},
{-32'd11899, 32'd5060, -32'd2692, -32'd12921},
{32'd1316, 32'd10555, 32'd7206, 32'd3546},
{-32'd2471, -32'd2678, 32'd1666, -32'd891},
{-32'd10300, -32'd2895, -32'd9445, -32'd3791},
{-32'd16485, -32'd10827, 32'd1464, -32'd9657},
{32'd9927, -32'd6488, -32'd4067, 32'd6652},
{32'd1858, 32'd9276, -32'd5082, 32'd5838},
{-32'd8011, 32'd6728, -32'd13473, 32'd5102},
{32'd7581, 32'd9119, 32'd6848, 32'd8330},
{32'd8656, 32'd3696, 32'd9580, 32'd8386},
{-32'd7136, 32'd1663, -32'd4881, -32'd2634},
{-32'd2007, -32'd6681, 32'd7889, 32'd4941},
{32'd1368, -32'd5059, 32'd2847, -32'd6196},
{-32'd8194, 32'd2543, -32'd10328, -32'd7728},
{-32'd3152, 32'd1341, 32'd9385, 32'd2164},
{-32'd1347, -32'd3572, -32'd15654, 32'd3324},
{-32'd6887, -32'd495, 32'd8215, 32'd11000},
{32'd6317, -32'd13348, -32'd2147, -32'd8672},
{-32'd5968, -32'd7922, 32'd7435, 32'd8833},
{-32'd2514, -32'd2138, -32'd12377, -32'd1625},
{32'd370, -32'd684, -32'd5606, 32'd12973},
{-32'd12117, 32'd1186, 32'd71, -32'd3055},
{32'd2162, 32'd8386, 32'd621, 32'd8766},
{-32'd112, 32'd604, -32'd3366, 32'd3476},
{-32'd2184, -32'd9003, 32'd6184, -32'd3646},
{-32'd8470, 32'd4640, 32'd4418, -32'd824},
{32'd8971, -32'd3111, -32'd7542, 32'd2834},
{-32'd2703, 32'd6680, 32'd6215, -32'd5178},
{32'd4794, -32'd12788, 32'd223, -32'd9108},
{-32'd756, -32'd2558, -32'd4594, -32'd79},
{32'd4989, -32'd2529, 32'd1908, -32'd9921},
{-32'd4510, -32'd6293, 32'd5, -32'd3583},
{32'd9441, -32'd7803, -32'd11748, 32'd992},
{-32'd1510, 32'd8608, 32'd7679, -32'd2488},
{32'd10609, 32'd3365, -32'd4496, 32'd6542},
{-32'd1501, -32'd7003, 32'd3825, -32'd4676},
{32'd11915, 32'd1759, -32'd534, 32'd2743},
{-32'd2791, 32'd4797, -32'd1006, 32'd3480},
{-32'd1168, -32'd11318, -32'd5712, -32'd4454},
{-32'd1078, -32'd7046, 32'd2019, -32'd3847},
{-32'd389, 32'd7666, -32'd9761, 32'd8455},
{-32'd322, -32'd3356, -32'd2315, 32'd3921},
{-32'd2473, -32'd11250, 32'd711, -32'd5302},
{-32'd1884, -32'd2041, 32'd2842, -32'd6006},
{-32'd13538, 32'd3133, -32'd1712, -32'd47},
{32'd17295, 32'd3160, 32'd6940, -32'd5011},
{32'd17665, -32'd3167, 32'd10246, -32'd3698},
{-32'd9740, -32'd8317, 32'd547, -32'd10960},
{-32'd2047, 32'd3958, -32'd5677, -32'd7733},
{32'd4381, -32'd2105, -32'd7817, 32'd14315},
{-32'd7975, 32'd2806, -32'd3835, 32'd11860},
{-32'd17859, -32'd3058, -32'd7580, 32'd2145},
{32'd1383, 32'd3286, 32'd1673, 32'd3667},
{32'd14904, 32'd8306, 32'd9269, -32'd10702},
{-32'd8521, -32'd5375, -32'd2814, 32'd831},
{-32'd5167, 32'd5553, -32'd14890, 32'd1480},
{-32'd11675, -32'd9091, -32'd2532, -32'd2462},
{-32'd1475, -32'd8190, -32'd2495, -32'd2901},
{32'd4173, -32'd16294, -32'd3347, 32'd2242},
{32'd9931, -32'd2186, -32'd4979, -32'd5760},
{-32'd687, -32'd5981, -32'd7037, 32'd1229},
{32'd2981, 32'd13570, 32'd10199, 32'd5473},
{32'd713, -32'd5678, -32'd2536, -32'd114},
{-32'd6479, 32'd1852, 32'd4578, -32'd6193},
{-32'd1595, -32'd1403, -32'd5812, 32'd47},
{-32'd3341, 32'd2338, 32'd2228, -32'd637},
{32'd1833, 32'd6417, 32'd7911, 32'd10977},
{32'd3222, -32'd4241, 32'd5067, 32'd3215},
{-32'd4008, -32'd6508, -32'd4921, 32'd7152},
{32'd2223, -32'd6400, -32'd8012, -32'd7598},
{-32'd7109, -32'd11334, -32'd5757, 32'd7133},
{32'd5629, 32'd7809, 32'd3697, -32'd2795},
{32'd5366, 32'd1760, 32'd2455, 32'd4272},
{32'd3488, -32'd748, -32'd5047, -32'd3174},
{-32'd2278, 32'd3186, -32'd8059, 32'd8127},
{-32'd5483, 32'd4693, 32'd6637, 32'd9084},
{-32'd4509, -32'd820, -32'd4193, 32'd8125},
{-32'd5198, 32'd3079, 32'd14218, 32'd5238},
{-32'd2411, -32'd6882, -32'd8421, -32'd1484},
{32'd907, 32'd3991, -32'd8195, 32'd5634},
{32'd9985, -32'd4671, 32'd421, -32'd3073},
{-32'd7590, -32'd1606, -32'd3242, -32'd4340},
{32'd4761, 32'd3649, 32'd1223, 32'd6766},
{32'd1743, -32'd7315, 32'd6553, 32'd5584},
{-32'd11330, -32'd1999, -32'd6981, -32'd1396},
{-32'd11106, 32'd6833, -32'd5506, 32'd1784},
{32'd3179, 32'd1284, 32'd8538, 32'd889},
{32'd3520, 32'd701, -32'd7470, 32'd6037},
{-32'd8914, 32'd2310, 32'd3419, -32'd7643},
{-32'd8842, -32'd7941, -32'd6577, 32'd2091},
{32'd4604, -32'd6700, -32'd15450, 32'd410},
{-32'd10831, -32'd7708, 32'd1949, 32'd4737},
{-32'd4542, -32'd5817, 32'd3051, 32'd9888},
{32'd5098, 32'd1207, 32'd5279, -32'd5122},
{-32'd299, -32'd4281, 32'd4039, 32'd6286},
{32'd8602, 32'd5719, -32'd2506, 32'd7158},
{-32'd1250, -32'd2632, 32'd5427, 32'd3779},
{32'd3352, 32'd6955, 32'd17080, 32'd3680},
{32'd1617, 32'd2973, -32'd4606, -32'd4781},
{-32'd2003, 32'd3082, 32'd4824, 32'd2261},
{32'd4703, 32'd376, -32'd1917, 32'd1990},
{32'd1958, 32'd6161, -32'd8402, 32'd3772},
{32'd5230, 32'd5667, -32'd551, -32'd1548},
{32'd1064, 32'd632, 32'd1840, -32'd9889},
{-32'd5739, -32'd14606, -32'd18707, -32'd1674},
{32'd8876, 32'd656, 32'd871, 32'd1666},
{-32'd7013, -32'd7072, -32'd5656, 32'd4246},
{-32'd86, -32'd2428, -32'd1641, 32'd9285},
{-32'd6430, 32'd2131, 32'd450, 32'd5085},
{32'd691, 32'd6572, 32'd1928, 32'd10764},
{-32'd6195, -32'd2182, 32'd3973, 32'd6162},
{32'd9140, 32'd7618, 32'd10510, -32'd2477},
{-32'd565, -32'd6804, -32'd1251, -32'd471},
{32'd6174, -32'd3043, -32'd6193, -32'd5658},
{32'd730, -32'd6909, 32'd6597, -32'd6847},
{32'd3203, 32'd1959, -32'd2234, -32'd2249},
{-32'd4809, -32'd5975, 32'd4742, -32'd2704},
{32'd12654, -32'd1980, 32'd4310, 32'd3969},
{-32'd2152, 32'd3186, 32'd1665, -32'd5961},
{-32'd5284, -32'd2625, -32'd9265, -32'd5803},
{-32'd11541, -32'd4472, 32'd5240, -32'd1540},
{32'd13781, 32'd5289, 32'd1703, 32'd6308},
{-32'd5432, -32'd122, -32'd15572, 32'd7449},
{32'd5170, 32'd5948, 32'd6972, 32'd6687},
{-32'd9836, -32'd4090, -32'd17282, 32'd295},
{32'd2025, 32'd73, 32'd3704, 32'd767},
{-32'd3875, 32'd2458, 32'd2895, 32'd4537},
{32'd2077, 32'd19089, -32'd2429, 32'd2699},
{-32'd1344, -32'd2056, 32'd4332, -32'd12845},
{-32'd5421, -32'd4977, 32'd1457, -32'd16793},
{-32'd12242, 32'd2214, 32'd4830, 32'd4832},
{-32'd8924, -32'd10577, -32'd3841, -32'd4190},
{32'd15480, 32'd3404, 32'd6247, 32'd3189},
{32'd9391, 32'd3307, 32'd3343, 32'd11162},
{-32'd14882, -32'd4742, -32'd1634, -32'd6376},
{32'd1181, -32'd11130, -32'd5157, -32'd4619},
{-32'd1802, -32'd1631, 32'd1939, -32'd4689},
{32'd6451, 32'd6872, -32'd2633, 32'd2976},
{32'd13092, 32'd658, 32'd11517, 32'd1570},
{-32'd3547, -32'd12633, -32'd3738, -32'd10287},
{-32'd6026, -32'd3548, -32'd1770, -32'd2988},
{-32'd2426, 32'd4083, -32'd3212, 32'd4759},
{32'd3592, -32'd14537, -32'd3681, 32'd1458},
{-32'd7360, -32'd13094, -32'd2666, -32'd9227},
{-32'd3065, -32'd1442, -32'd1432, 32'd1399},
{-32'd6318, -32'd7262, -32'd10382, -32'd10747},
{32'd3156, 32'd8451, 32'd7680, 32'd9017},
{-32'd4750, -32'd3103, -32'd5014, -32'd8329},
{32'd646, 32'd5169, -32'd4873, 32'd3387},
{-32'd558, 32'd2284, -32'd8844, 32'd1578},
{-32'd7280, -32'd2905, -32'd6657, -32'd646},
{-32'd1480, 32'd3548, -32'd675, -32'd7106},
{32'd8730, 32'd9175, 32'd105, -32'd4788},
{-32'd6321, 32'd7556, 32'd3078, 32'd4497},
{32'd3556, 32'd9671, -32'd1249, -32'd4158},
{-32'd1501, 32'd6181, -32'd1453, 32'd863},
{-32'd5977, -32'd7032, 32'd11555, 32'd3485},
{-32'd1205, -32'd270, -32'd3989, -32'd7192},
{-32'd5739, 32'd3483, -32'd7966, -32'd3830},
{32'd15015, -32'd5322, 32'd7061, 32'd12246},
{-32'd3661, 32'd7022, 32'd9151, 32'd3044},
{-32'd145, -32'd2505, 32'd3231, 32'd1871},
{-32'd1562, 32'd4817, -32'd7308, -32'd664},
{32'd6851, -32'd4899, -32'd15262, -32'd4019},
{32'd3132, -32'd6430, -32'd4028, -32'd328},
{32'd7045, 32'd12766, 32'd8575, 32'd7596},
{32'd2134, 32'd5432, -32'd5152, -32'd1918},
{-32'd3430, -32'd2886, -32'd6427, -32'd7062},
{32'd5108, -32'd4095, -32'd7925, -32'd565},
{-32'd616, 32'd15712, 32'd3539, -32'd5057},
{32'd9884, 32'd3962, -32'd1641, 32'd8093},
{32'd12552, -32'd3114, 32'd10631, 32'd920},
{32'd13364, -32'd346, 32'd5954, 32'd4895},
{32'd1597, 32'd445, 32'd1217, 32'd8385},
{-32'd1529, -32'd11643, -32'd6081, -32'd8291},
{32'd2178, -32'd3550, -32'd1278, 32'd7608},
{32'd4776, -32'd5768, -32'd12905, -32'd11662},
{-32'd9113, 32'd576, 32'd3614, -32'd2180},
{32'd1622, -32'd5308, -32'd9453, 32'd3682},
{-32'd5292, 32'd5039, 32'd2695, 32'd362},
{32'd8871, 32'd5406, 32'd2827, 32'd1041},
{-32'd2278, -32'd593, -32'd3671, -32'd1919},
{-32'd10770, 32'd1489, -32'd4479, 32'd3065},
{-32'd860, -32'd7864, 32'd4255, 32'd1150},
{-32'd3174, -32'd6331, 32'd4785, -32'd1886},
{-32'd9700, -32'd7618, -32'd8988, -32'd12297},
{-32'd12184, 32'd12579, 32'd3119, -32'd4699},
{32'd9720, -32'd998, -32'd3107, 32'd3225},
{-32'd7987, -32'd108, -32'd13408, -32'd2513}
},
{{32'd5794, -32'd982, 32'd4654, -32'd7126},
{-32'd3796, -32'd9415, 32'd4407, -32'd8974},
{32'd8431, 32'd534, -32'd9680, -32'd6215},
{32'd4229, -32'd2727, -32'd3656, -32'd3494},
{-32'd6536, 32'd4204, 32'd16438, 32'd224},
{32'd6380, -32'd4854, 32'd1053, -32'd7576},
{32'd8555, 32'd8359, 32'd4551, -32'd5061},
{-32'd5605, -32'd4813, -32'd2112, -32'd7908},
{32'd10263, -32'd1365, -32'd5778, -32'd6338},
{32'd10533, -32'd3861, 32'd1430, -32'd28},
{-32'd8892, 32'd10054, -32'd2259, -32'd538},
{32'd3913, -32'd2155, -32'd1292, 32'd5418},
{32'd1792, -32'd3360, 32'd16690, -32'd4569},
{32'd2998, 32'd6828, -32'd2337, 32'd1671},
{-32'd13099, 32'd5047, -32'd5498, 32'd14156},
{-32'd15689, 32'd8057, 32'd4030, 32'd5017},
{32'd7796, 32'd10488, 32'd4946, -32'd6548},
{32'd5836, -32'd7945, -32'd8032, 32'd5267},
{-32'd8001, 32'd6614, 32'd3361, -32'd4913},
{32'd4455, 32'd2446, -32'd1643, -32'd9918},
{32'd6246, 32'd6707, 32'd16517, -32'd10879},
{-32'd8561, 32'd7352, 32'd2174, -32'd5357},
{-32'd11874, -32'd1761, 32'd5789, -32'd2713},
{-32'd6694, -32'd2416, -32'd10796, 32'd2615},
{32'd3992, -32'd6117, 32'd3977, -32'd8122},
{32'd1090, 32'd6309, 32'd4039, -32'd4947},
{-32'd8898, -32'd11571, -32'd1571, 32'd1807},
{32'd1875, 32'd2797, 32'd8674, 32'd7558},
{32'd3973, 32'd6118, 32'd23243, 32'd2686},
{-32'd1129, 32'd9821, 32'd2761, 32'd2343},
{-32'd6501, 32'd13518, 32'd10059, -32'd951},
{32'd1816, 32'd2194, 32'd5894, -32'd5862},
{32'd5026, 32'd2989, -32'd3537, 32'd3308},
{-32'd1409, 32'd808, -32'd8401, 32'd11526},
{32'd13194, -32'd1586, 32'd6401, 32'd2941},
{32'd7821, 32'd880, 32'd6843, -32'd11114},
{-32'd5731, 32'd8349, 32'd7272, -32'd6012},
{32'd8742, 32'd5026, -32'd5229, -32'd4483},
{-32'd740, 32'd8770, -32'd3358, -32'd6018},
{-32'd6224, -32'd3813, 32'd2528, 32'd1408},
{-32'd13476, 32'd70, -32'd6657, -32'd158},
{32'd2198, -32'd514, -32'd3659, 32'd4046},
{-32'd2524, -32'd6158, -32'd2731, -32'd8498},
{-32'd2608, -32'd936, 32'd3484, 32'd1781},
{32'd1222, -32'd17910, -32'd8577, 32'd4067},
{-32'd5076, 32'd2841, 32'd2506, 32'd1076},
{32'd1546, -32'd4001, 32'd2723, 32'd1952},
{-32'd6018, -32'd7692, -32'd4918, 32'd5005},
{32'd2499, -32'd4960, -32'd4038, -32'd13440},
{-32'd5959, -32'd2772, 32'd4825, -32'd10067},
{32'd1537, 32'd218, -32'd5146, -32'd2284},
{-32'd4138, -32'd2550, -32'd8176, 32'd1484},
{-32'd3965, -32'd2635, -32'd1904, 32'd13453},
{32'd2760, -32'd2659, -32'd5290, -32'd6321},
{32'd2128, -32'd6215, 32'd6723, 32'd16455},
{-32'd408, 32'd10220, 32'd3718, -32'd11391},
{32'd5365, 32'd10471, -32'd4160, -32'd1567},
{-32'd2449, 32'd9852, -32'd8720, -32'd3234},
{-32'd9798, 32'd6164, -32'd15126, -32'd3569},
{-32'd10641, -32'd3069, 32'd7402, -32'd6535},
{-32'd8317, -32'd6795, 32'd11048, 32'd9108},
{-32'd7518, 32'd2614, -32'd889, 32'd5942},
{-32'd6227, 32'd2755, 32'd386, -32'd4450},
{-32'd2865, -32'd4601, 32'd10617, -32'd6499},
{-32'd1887, 32'd1843, -32'd5576, -32'd740},
{32'd7980, -32'd2072, 32'd966, 32'd9288},
{-32'd11783, 32'd6187, 32'd4029, 32'd8235},
{-32'd9192, -32'd8998, -32'd6805, 32'd13774},
{-32'd5128, -32'd12622, -32'd7114, 32'd3724},
{32'd3668, 32'd369, 32'd8565, 32'd9421},
{-32'd6979, -32'd842, 32'd1834, 32'd10265},
{32'd1935, 32'd6341, -32'd5829, 32'd10214},
{-32'd4762, 32'd7817, -32'd8115, -32'd1991},
{-32'd6762, 32'd12313, 32'd2408, -32'd1806},
{32'd4231, -32'd2717, -32'd1108, 32'd3993},
{-32'd6981, 32'd302, -32'd3146, 32'd6099},
{-32'd7662, 32'd6300, -32'd7232, -32'd7651},
{-32'd12244, 32'd1719, 32'd14179, -32'd7757},
{-32'd2612, 32'd3046, 32'd2466, -32'd4614},
{-32'd2150, -32'd5011, -32'd1571, -32'd2881},
{-32'd1452, -32'd10394, -32'd8074, 32'd1268},
{32'd1609, -32'd6355, 32'd4578, -32'd17689},
{-32'd802, 32'd12081, 32'd12450, -32'd1731},
{32'd4202, 32'd2230, -32'd8215, 32'd7224},
{-32'd59, 32'd363, -32'd517, -32'd1348},
{32'd2648, 32'd4571, -32'd2234, 32'd8954},
{32'd9186, -32'd12116, -32'd8738, -32'd10129},
{-32'd13908, 32'd6164, 32'd2888, -32'd3879},
{-32'd3842, 32'd3138, -32'd7440, -32'd1006},
{-32'd12110, -32'd7437, 32'd6895, 32'd4467},
{32'd4559, 32'd1653, -32'd6156, -32'd5377},
{-32'd189, 32'd9980, -32'd1213, -32'd7794},
{-32'd2223, -32'd5614, 32'd1769, 32'd5777},
{32'd10047, -32'd1991, -32'd5277, 32'd8074},
{32'd44, 32'd247, 32'd9962, 32'd13117},
{-32'd15517, -32'd8782, -32'd11655, -32'd5358},
{32'd6736, 32'd2873, -32'd5404, -32'd6306},
{32'd11945, -32'd5271, 32'd9930, -32'd3856},
{-32'd2945, 32'd8253, 32'd18125, 32'd7710},
{32'd3855, -32'd4491, 32'd35, 32'd1891},
{-32'd9617, -32'd3590, -32'd4381, -32'd6090},
{32'd9281, 32'd719, 32'd3277, 32'd11980},
{32'd9948, 32'd294, -32'd2179, 32'd6126},
{-32'd6131, -32'd3899, 32'd2344, -32'd565},
{-32'd11207, 32'd9075, -32'd2444, -32'd1780},
{-32'd5831, -32'd7909, -32'd3244, 32'd4698},
{32'd9278, 32'd5792, 32'd6568, -32'd8493},
{32'd3741, 32'd2622, 32'd1450, 32'd3003},
{32'd2689, -32'd10418, 32'd6160, 32'd2358},
{-32'd4100, 32'd3000, 32'd2478, 32'd3052},
{-32'd14831, -32'd49, -32'd5712, 32'd4773},
{-32'd678, 32'd508, -32'd3601, -32'd10398},
{32'd10434, -32'd485, -32'd3098, -32'd3579},
{32'd8665, -32'd2895, -32'd2530, 32'd502},
{-32'd3559, -32'd5152, 32'd2807, -32'd3074},
{-32'd9975, 32'd2132, 32'd3978, 32'd3798},
{32'd7699, 32'd7433, 32'd7059, 32'd1333},
{32'd8347, -32'd9326, 32'd3610, 32'd1373},
{32'd1461, 32'd10795, 32'd7837, 32'd7257},
{32'd5041, 32'd7097, 32'd5179, 32'd6573},
{32'd572, -32'd757, 32'd1711, -32'd1237},
{32'd923, 32'd6202, -32'd7286, 32'd8599},
{-32'd2909, -32'd12, 32'd5062, 32'd2944},
{32'd509, 32'd5710, 32'd4415, -32'd5616},
{-32'd6139, -32'd3448, 32'd1102, -32'd10627},
{32'd3862, -32'd8666, -32'd4946, -32'd797},
{-32'd5696, 32'd498, 32'd2754, -32'd12319},
{32'd2143, -32'd1334, -32'd4922, -32'd2213},
{-32'd7766, -32'd7716, 32'd2081, -32'd1004},
{32'd3247, -32'd5077, 32'd52, -32'd2015},
{-32'd7447, 32'd940, 32'd17381, -32'd302},
{32'd7196, -32'd3214, 32'd4512, 32'd4338},
{-32'd9116, -32'd1243, -32'd1873, -32'd4692},
{-32'd6340, 32'd3475, 32'd3788, -32'd737},
{-32'd929, -32'd7492, -32'd1548, 32'd6732},
{32'd5020, 32'd2722, -32'd407, 32'd1654},
{32'd2679, -32'd251, 32'd4410, -32'd504},
{32'd12749, -32'd15712, 32'd4371, -32'd8743},
{32'd3323, 32'd3308, -32'd7073, 32'd2452},
{-32'd19279, -32'd5336, 32'd244, -32'd6961},
{-32'd8522, -32'd15107, -32'd5639, -32'd2102},
{-32'd3954, 32'd8849, -32'd1477, -32'd9129},
{-32'd3018, 32'd4963, 32'd3362, 32'd4203},
{-32'd11988, 32'd4476, 32'd12856, 32'd2595},
{32'd5532, -32'd217, 32'd6973, -32'd3287},
{-32'd8821, 32'd3890, -32'd9765, 32'd2342},
{-32'd6271, -32'd20, -32'd10385, -32'd7393},
{-32'd3421, 32'd5301, 32'd4312, -32'd1116},
{32'd5139, 32'd3943, 32'd9627, -32'd595},
{32'd740, -32'd9210, 32'd5225, -32'd14669},
{-32'd5555, -32'd1837, -32'd7944, 32'd1480},
{32'd11720, -32'd2825, -32'd1879, -32'd1294},
{32'd1251, 32'd5932, -32'd2667, -32'd887},
{-32'd2061, -32'd3068, -32'd4439, -32'd1289},
{-32'd4701, -32'd5360, -32'd8350, 32'd1569},
{-32'd3502, -32'd2088, -32'd1321, 32'd7686},
{32'd8973, 32'd1103, 32'd12803, -32'd8132},
{32'd13813, 32'd6477, -32'd8656, -32'd3271},
{-32'd411, -32'd5106, -32'd3955, -32'd6986},
{32'd4764, -32'd6102, 32'd7846, -32'd8668},
{32'd3877, 32'd3980, -32'd7853, -32'd7795},
{32'd1123, -32'd15189, 32'd4282, 32'd7613},
{-32'd5054, 32'd6019, 32'd13130, -32'd9819},
{32'd13066, -32'd2763, -32'd2833, -32'd1861},
{32'd4187, 32'd5696, 32'd20216, 32'd3791},
{-32'd472, 32'd3079, -32'd3272, -32'd743},
{-32'd2580, -32'd1309, 32'd9312, 32'd9351},
{-32'd6164, 32'd1522, -32'd1835, 32'd5132},
{-32'd1979, 32'd162, 32'd7394, 32'd1000},
{-32'd10129, 32'd9779, 32'd2060, 32'd10436},
{-32'd2575, 32'd5856, 32'd874, -32'd7911},
{32'd3448, -32'd4703, -32'd1444, -32'd15879},
{32'd15039, -32'd1597, 32'd8020, 32'd6523},
{-32'd6194, -32'd5463, -32'd17617, 32'd6003},
{32'd1607, -32'd4491, 32'd9962, -32'd9568},
{32'd4833, 32'd4793, -32'd1802, 32'd3059},
{32'd558, -32'd13394, -32'd171, 32'd4874},
{32'd5811, -32'd1826, 32'd12127, -32'd6273},
{32'd8490, -32'd2034, 32'd15083, 32'd5815},
{-32'd17001, 32'd4582, -32'd17755, 32'd7458},
{-32'd4104, -32'd10352, 32'd11458, -32'd11727},
{-32'd4191, 32'd1856, -32'd3185, -32'd2058},
{-32'd13885, -32'd5797, 32'd8337, -32'd8720},
{-32'd10591, -32'd15844, -32'd657, 32'd730},
{-32'd5837, -32'd7593, -32'd8858, 32'd5923},
{32'd7504, 32'd2804, 32'd2787, 32'd5050},
{32'd14236, -32'd1734, 32'd14971, 32'd3565},
{32'd7838, 32'd4105, 32'd6327, 32'd2033},
{-32'd319, 32'd17635, 32'd8191, -32'd6581},
{32'd849, 32'd15586, 32'd2187, -32'd6054},
{-32'd966, 32'd10482, -32'd5073, -32'd10885},
{32'd1552, 32'd6190, -32'd4867, -32'd1413},
{-32'd10802, -32'd100, -32'd13017, 32'd13118},
{-32'd7529, -32'd3026, 32'd9723, -32'd11461},
{32'd834, -32'd10601, -32'd4370, 32'd7522},
{32'd4083, -32'd10722, -32'd4790, -32'd7308},
{-32'd1122, -32'd5763, -32'd3360, -32'd6151},
{-32'd8197, 32'd303, 32'd997, 32'd13196},
{-32'd8957, 32'd12693, -32'd1548, -32'd2335},
{-32'd300, -32'd13465, -32'd12174, -32'd3170},
{-32'd8337, -32'd389, -32'd5609, -32'd4299},
{-32'd2431, 32'd2882, -32'd3286, 32'd4887},
{32'd3502, -32'd4608, 32'd1287, 32'd4331},
{32'd12532, 32'd5893, -32'd516, 32'd2919},
{-32'd3679, 32'd1240, -32'd11473, 32'd3934},
{32'd6083, 32'd3548, 32'd4264, 32'd4721},
{-32'd1610, 32'd5978, 32'd4588, -32'd4596},
{-32'd7896, 32'd6030, -32'd7796, 32'd3147},
{32'd6828, 32'd6645, 32'd2275, 32'd2075},
{32'd1865, -32'd10769, 32'd3332, 32'd7438},
{-32'd3365, 32'd2477, -32'd18920, -32'd2539},
{32'd5055, -32'd4056, 32'd833, -32'd1639},
{32'd7070, 32'd3324, 32'd4119, -32'd7821},
{32'd7664, -32'd5560, -32'd10871, 32'd6267},
{-32'd11848, -32'd10178, -32'd11481, -32'd7168},
{-32'd380, -32'd898, -32'd2889, -32'd2643},
{32'd9716, 32'd1063, -32'd4413, 32'd4707},
{-32'd12242, 32'd5444, 32'd5562, 32'd7158},
{32'd9683, 32'd4094, 32'd5521, 32'd440},
{32'd239, -32'd7865, -32'd2054, 32'd19234},
{32'd2231, 32'd9089, -32'd13077, 32'd3702},
{32'd2938, -32'd2365, 32'd3144, 32'd1822},
{32'd8268, 32'd5886, 32'd11776, -32'd2749},
{32'd6235, 32'd10139, 32'd2988, 32'd2192},
{-32'd1637, 32'd13862, 32'd12142, 32'd550},
{32'd3564, -32'd7981, -32'd615, -32'd703},
{-32'd7039, 32'd1381, -32'd3504, 32'd7985},
{-32'd3841, -32'd13199, -32'd1893, -32'd4566},
{32'd6917, -32'd9983, -32'd12486, 32'd11705},
{-32'd4162, 32'd574, -32'd1193, 32'd8817},
{-32'd2771, 32'd6212, 32'd2488, -32'd98},
{-32'd1107, 32'd11725, -32'd2911, 32'd6492},
{-32'd5608, 32'd7890, 32'd5104, -32'd9039},
{32'd11430, 32'd591, -32'd6249, 32'd4829},
{32'd11315, -32'd10182, -32'd9184, 32'd169},
{-32'd8524, -32'd7055, -32'd13915, 32'd5929},
{32'd5440, -32'd4156, -32'd3904, 32'd2048},
{32'd905, 32'd8314, 32'd5391, -32'd4243},
{32'd1096, 32'd7189, 32'd6095, 32'd8103},
{32'd1537, 32'd11082, 32'd4686, 32'd4260},
{-32'd2961, 32'd339, 32'd7574, 32'd2134},
{32'd155, 32'd2004, -32'd6286, 32'd3967},
{-32'd17094, 32'd399, -32'd484, 32'd2664},
{-32'd6312, 32'd16936, -32'd10992, 32'd2222},
{32'd10373, 32'd2263, 32'd11149, 32'd3399},
{-32'd16495, 32'd595, -32'd950, 32'd5293},
{-32'd3879, 32'd4003, -32'd9627, -32'd7219},
{32'd959, -32'd6488, -32'd7522, -32'd7998},
{32'd3856, 32'd2773, 32'd2242, 32'd3851},
{-32'd4499, 32'd7873, 32'd1617, 32'd5135},
{-32'd6669, -32'd1843, -32'd6042, -32'd5525},
{32'd6881, -32'd5377, 32'd2381, -32'd9824},
{32'd670, -32'd4137, -32'd8580, 32'd3092},
{-32'd6948, 32'd7054, -32'd1316, -32'd4867},
{-32'd6575, 32'd12565, -32'd523, 32'd2600},
{32'd18559, 32'd462, 32'd6052, -32'd458},
{-32'd5592, -32'd9647, -32'd5606, 32'd2681},
{32'd5106, 32'd677, 32'd8433, 32'd2353},
{-32'd1623, 32'd1419, -32'd16762, -32'd5535},
{32'd7721, -32'd2701, -32'd5913, 32'd7946},
{32'd21587, 32'd2107, 32'd9263, -32'd2594},
{32'd9615, 32'd1516, 32'd3039, 32'd4755},
{-32'd3904, -32'd13743, -32'd1808, -32'd6545},
{-32'd17401, -32'd12256, -32'd6196, 32'd3092},
{32'd6842, 32'd4803, -32'd1494, -32'd476},
{32'd9606, -32'd2657, 32'd3418, -32'd17446},
{32'd7378, -32'd1382, -32'd241, -32'd4215},
{32'd2238, 32'd9858, 32'd2064, 32'd2703},
{32'd5943, 32'd994, -32'd7827, 32'd8575},
{32'd484, 32'd1199, -32'd6285, 32'd1620},
{32'd2452, 32'd10947, -32'd3688, 32'd20819},
{32'd1992, -32'd1546, -32'd6730, 32'd10955},
{-32'd5817, -32'd3644, 32'd5525, -32'd129},
{-32'd5924, 32'd7754, 32'd5664, 32'd2029},
{-32'd6326, 32'd17285, -32'd16498, -32'd1925},
{-32'd3771, 32'd14714, -32'd714, 32'd939},
{32'd11553, -32'd955, 32'd4571, -32'd1504},
{-32'd4986, 32'd10085, 32'd7484, 32'd7518},
{-32'd11510, -32'd1622, -32'd2814, 32'd788},
{-32'd9233, -32'd7091, 32'd8358, -32'd382},
{32'd5607, -32'd7911, 32'd11492, -32'd5348},
{-32'd4615, 32'd6748, 32'd3745, -32'd9339},
{-32'd3222, 32'd15049, 32'd3869, 32'd1274},
{-32'd10459, 32'd380, 32'd3286, 32'd2811},
{32'd2043, 32'd8817, 32'd7251, 32'd6820},
{-32'd9936, -32'd2926, -32'd14739, -32'd3093},
{32'd7363, -32'd4990, -32'd4110, -32'd2165},
{-32'd9140, -32'd978, -32'd9471, -32'd2462},
{32'd364, 32'd720, -32'd8281, -32'd7655},
{-32'd3957, 32'd6190, -32'd10566, 32'd4165},
{32'd4977, 32'd4405, 32'd3221, 32'd1027},
{-32'd49, -32'd7260, 32'd1312, -32'd10892},
{-32'd1094, 32'd7220, -32'd1869, -32'd17077},
{32'd3495, -32'd5968, -32'd2396, -32'd7814},
{-32'd5994, 32'd8610, -32'd3367, 32'd9904},
{-32'd4939, 32'd4690, -32'd11482, 32'd7388},
{32'd525, -32'd2454, -32'd13456, -32'd8763},
{32'd13217, -32'd5282, 32'd1474, -32'd3311},
{32'd2851, -32'd5038, 32'd13506, 32'd7422},
{-32'd12045, 32'd7351, -32'd409, -32'd12154}
},
{{-32'd5321, -32'd5665, 32'd4281, 32'd8100},
{32'd9859, 32'd3549, 32'd2409, -32'd3781},
{-32'd4450, -32'd2641, 32'd3752, -32'd4592},
{32'd13280, 32'd14836, 32'd8378, 32'd8262},
{-32'd512, 32'd12864, 32'd4472, -32'd3631},
{-32'd3239, -32'd7193, -32'd3106, 32'd1755},
{32'd4273, 32'd8327, 32'd6252, 32'd2658},
{32'd2702, -32'd1261, -32'd460, -32'd5586},
{32'd1400, -32'd10136, 32'd7300, 32'd8708},
{32'd14098, 32'd7517, 32'd12565, 32'd3475},
{32'd2468, 32'd2669, -32'd11286, -32'd2077},
{-32'd9952, -32'd2875, -32'd514, -32'd6412},
{-32'd11370, 32'd9735, 32'd5544, -32'd130},
{32'd4659, -32'd716, 32'd838, -32'd11338},
{-32'd7944, 32'd9384, -32'd8301, 32'd4042},
{-32'd5333, 32'd3253, 32'd92, 32'd6999},
{32'd140, -32'd9670, 32'd10629, 32'd4329},
{32'd2069, -32'd5208, 32'd2278, 32'd1235},
{-32'd4330, 32'd4494, -32'd10701, -32'd13843},
{-32'd6964, 32'd6176, -32'd11401, 32'd1158},
{-32'd3933, -32'd1296, -32'd7842, -32'd3569},
{32'd4979, 32'd1017, -32'd8377, 32'd5687},
{32'd845, 32'd5429, 32'd4266, 32'd5791},
{-32'd6344, -32'd464, -32'd11491, 32'd535},
{32'd1530, 32'd915, 32'd1190, 32'd8130},
{-32'd4125, 32'd8199, -32'd7326, -32'd2174},
{32'd2651, -32'd16362, -32'd878, 32'd3999},
{-32'd1519, 32'd11587, 32'd7489, 32'd7327},
{32'd7776, 32'd5869, 32'd6375, -32'd1738},
{-32'd457, 32'd4769, -32'd1133, -32'd343},
{-32'd8207, 32'd10868, -32'd544, -32'd5851},
{-32'd5190, 32'd2060, -32'd10250, 32'd1167},
{-32'd2758, 32'd12914, 32'd3783, -32'd4961},
{-32'd11990, 32'd831, -32'd11510, -32'd5887},
{32'd981, 32'd7718, 32'd14584, 32'd4880},
{32'd1906, -32'd8497, -32'd5871, 32'd1421},
{-32'd6187, 32'd7325, 32'd6152, 32'd2712},
{32'd7780, -32'd5038, -32'd5741, -32'd1922},
{-32'd2164, 32'd8682, 32'd5593, 32'd2244},
{-32'd5371, -32'd6913, 32'd4059, 32'd6165},
{32'd8074, -32'd2620, -32'd2977, -32'd310},
{32'd4738, 32'd3535, -32'd3234, 32'd192},
{32'd5754, -32'd12044, 32'd4602, 32'd4433},
{-32'd6291, -32'd11025, -32'd3560, 32'd1435},
{-32'd7781, -32'd2178, -32'd7328, -32'd14707},
{32'd2912, 32'd4578, -32'd9169, -32'd2604},
{-32'd2485, 32'd1745, -32'd7627, -32'd4071},
{-32'd19391, -32'd6460, 32'd3188, -32'd7582},
{32'd3451, 32'd5948, 32'd12037, 32'd2951},
{-32'd1547, -32'd1285, -32'd3005, -32'd123},
{32'd172, -32'd8691, -32'd2339, -32'd1850},
{32'd4638, 32'd4465, -32'd10037, 32'd7245},
{-32'd6201, 32'd2546, -32'd4860, -32'd5170},
{32'd6069, 32'd2079, 32'd5697, 32'd522},
{32'd1148, 32'd7042, 32'd8968, 32'd4654},
{32'd7997, 32'd2243, -32'd5507, -32'd5296},
{-32'd8952, -32'd421, 32'd12526, 32'd3577},
{-32'd5268, 32'd6283, -32'd9238, 32'd800},
{32'd3157, 32'd6993, -32'd4983, -32'd4794},
{-32'd5331, -32'd7977, 32'd2564, -32'd1696},
{-32'd1366, 32'd1152, -32'd3687, 32'd74},
{32'd10425, 32'd5170, 32'd14247, 32'd733},
{32'd1565, -32'd5264, -32'd2849, -32'd4129},
{32'd6197, 32'd6661, -32'd4593, 32'd2994},
{-32'd9120, 32'd861, 32'd1332, 32'd2163},
{32'd943, 32'd1924, 32'd10093, 32'd11583},
{-32'd10086, -32'd1608, -32'd9332, 32'd3435},
{-32'd11218, -32'd7144, -32'd226, 32'd1857},
{-32'd8233, -32'd1430, -32'd6020, -32'd10094},
{32'd17627, -32'd3491, 32'd3981, -32'd4375},
{-32'd11872, 32'd11437, -32'd8637, -32'd565},
{32'd4699, 32'd3072, 32'd738, 32'd940},
{-32'd4539, 32'd1065, -32'd10252, -32'd4374},
{-32'd4981, 32'd386, 32'd2310, 32'd9738},
{32'd6666, -32'd802, 32'd4070, 32'd8167},
{-32'd4094, -32'd6448, 32'd2236, 32'd6454},
{32'd4603, -32'd3469, -32'd5068, -32'd5333},
{-32'd14815, 32'd10549, -32'd9825, -32'd1465},
{32'd10070, 32'd3423, 32'd13161, 32'd7751},
{-32'd328, -32'd7910, 32'd729, -32'd6817},
{32'd1326, -32'd196, 32'd7513, 32'd8343},
{-32'd1717, -32'd2589, 32'd7160, 32'd7781},
{-32'd2323, -32'd2591, -32'd9632, -32'd4935},
{-32'd498, -32'd2408, 32'd4639, -32'd2853},
{-32'd2568, -32'd8084, -32'd2445, -32'd7355},
{-32'd7530, 32'd205, -32'd10830, -32'd8921},
{-32'd2965, 32'd10880, 32'd2569, 32'd6014},
{-32'd10508, 32'd4153, -32'd11291, -32'd2995},
{32'd2498, 32'd1983, -32'd10156, -32'd8407},
{-32'd4650, -32'd8528, 32'd4849, -32'd11409},
{32'd6052, 32'd8200, 32'd3220, 32'd6675},
{32'd10316, -32'd1333, -32'd6406, 32'd7102},
{-32'd1947, 32'd2368, 32'd473, -32'd11835},
{32'd2511, 32'd4778, 32'd14667, 32'd2228},
{32'd589, 32'd8137, 32'd6569, -32'd4416},
{-32'd4916, 32'd7484, -32'd3532, -32'd2066},
{32'd3021, 32'd13935, 32'd680, -32'd306},
{32'd8619, -32'd10989, 32'd804, -32'd1376},
{-32'd11477, 32'd11201, 32'd5543, -32'd1029},
{32'd8610, 32'd5744, 32'd8812, -32'd954},
{32'd1216, -32'd4270, -32'd8363, -32'd3022},
{32'd2359, -32'd16899, 32'd1636, -32'd1912},
{32'd227, -32'd4289, 32'd132, 32'd6221},
{32'd3014, -32'd4269, 32'd2683, 32'd10331},
{32'd4110, 32'd2119, -32'd3921, -32'd2087},
{-32'd5909, 32'd7761, -32'd2017, 32'd4092},
{32'd3839, -32'd6123, 32'd6463, -32'd3232},
{-32'd5979, -32'd1598, 32'd3903, -32'd8019},
{32'd4595, 32'd2335, 32'd1844, 32'd2858},
{-32'd4533, -32'd7767, 32'd1112, -32'd13517},
{-32'd2593, 32'd8589, 32'd3579, 32'd861},
{32'd623, -32'd2740, -32'd30, 32'd5276},
{-32'd6761, 32'd2800, 32'd3556, 32'd7874},
{-32'd4372, 32'd11448, -32'd3648, 32'd15112},
{32'd6376, -32'd4368, -32'd3925, -32'd13939},
{32'd3784, -32'd6461, 32'd7459, -32'd2402},
{32'd4431, -32'd303, 32'd1136, -32'd2297},
{32'd1384, -32'd5331, 32'd3027, 32'd4907},
{32'd12386, -32'd9411, 32'd6914, 32'd5368},
{32'd6229, -32'd1691, 32'd13090, 32'd6656},
{-32'd18268, 32'd10970, 32'd2551, 32'd7970},
{32'd3296, 32'd5071, -32'd3011, -32'd1045},
{-32'd14788, -32'd5249, 32'd3808, -32'd263},
{32'd2772, -32'd6023, 32'd8718, -32'd9250},
{-32'd16572, -32'd315, -32'd6143, -32'd2329},
{32'd10214, 32'd6376, 32'd14469, 32'd17348},
{32'd653, -32'd16021, 32'd13, -32'd3582},
{-32'd5942, -32'd3920, -32'd10418, -32'd5199},
{-32'd3224, 32'd949, -32'd8370, 32'd4829},
{32'd2188, 32'd4688, -32'd9283, -32'd1732},
{-32'd2798, 32'd978, -32'd1670, -32'd846},
{-32'd14011, 32'd3513, -32'd8797, -32'd12638},
{-32'd607, -32'd5406, -32'd3504, -32'd3210},
{32'd12546, -32'd5350, 32'd8005, 32'd4441},
{-32'd3115, 32'd8408, -32'd1534, 32'd3200},
{32'd4602, -32'd2953, 32'd3972, -32'd11942},
{32'd1322, 32'd15582, -32'd3450, -32'd7785},
{-32'd8399, 32'd474, -32'd11695, 32'd871},
{32'd868, -32'd5551, 32'd8663, -32'd325},
{-32'd1196, 32'd1877, -32'd3737, -32'd4759},
{-32'd6170, 32'd2701, -32'd7535, -32'd2036},
{32'd8641, -32'd3272, 32'd677, -32'd10502},
{-32'd4915, 32'd5082, 32'd4402, 32'd7966},
{-32'd7945, 32'd307, -32'd18, 32'd10674},
{32'd10927, -32'd3000, 32'd9084, 32'd596},
{-32'd5433, 32'd7994, 32'd12428, 32'd12342},
{-32'd6190, 32'd4935, -32'd1333, -32'd10067},
{32'd9528, -32'd10202, 32'd3035, -32'd550},
{-32'd1958, -32'd15018, 32'd12959, 32'd7017},
{-32'd6319, -32'd10023, -32'd5912, -32'd6656},
{-32'd9851, 32'd2181, -32'd12871, -32'd1391},
{32'd9769, 32'd896, 32'd8226, 32'd7055},
{-32'd4855, -32'd10136, 32'd9349, -32'd78},
{32'd8940, 32'd3579, -32'd5524, -32'd4150},
{-32'd13688, 32'd4287, -32'd9890, -32'd1906},
{-32'd450, 32'd5287, 32'd4656, 32'd4493},
{-32'd2979, 32'd6073, -32'd7024, -32'd109},
{-32'd2590, -32'd282, -32'd2526, 32'd203},
{32'd1162, -32'd1328, 32'd7089, 32'd10857},
{-32'd737, 32'd15593, 32'd2042, -32'd3033},
{32'd2694, 32'd3739, -32'd129, -32'd3974},
{32'd5203, -32'd3060, 32'd7620, 32'd5090},
{32'd5823, -32'd897, -32'd2504, -32'd5734},
{32'd10919, 32'd744, 32'd12823, 32'd3905},
{32'd10893, -32'd5564, 32'd9046, 32'd4469},
{-32'd8459, -32'd11564, -32'd3176, 32'd5425},
{32'd5547, -32'd2947, 32'd15944, -32'd3868},
{-32'd4160, 32'd1805, -32'd5220, -32'd9012},
{-32'd4043, 32'd16082, -32'd3468, -32'd4431},
{32'd2553, -32'd10692, -32'd5052, 32'd3633},
{-32'd4507, -32'd2084, 32'd2776, 32'd5563},
{-32'd3763, -32'd5646, 32'd1850, -32'd6610},
{32'd2426, 32'd5172, 32'd10747, 32'd2678},
{32'd6655, -32'd7172, 32'd1996, -32'd1894},
{32'd17826, 32'd2156, -32'd4478, 32'd3208},
{-32'd10500, 32'd3617, 32'd1718, -32'd13276},
{32'd6091, -32'd7283, 32'd2793, -32'd3697},
{-32'd2078, 32'd939, 32'd8773, 32'd2968},
{32'd2975, -32'd9911, 32'd6264, 32'd6766},
{-32'd3533, 32'd2571, -32'd5069, 32'd1624},
{32'd6499, -32'd1562, 32'd649, 32'd1343},
{-32'd14605, 32'd10850, 32'd6086, 32'd810},
{-32'd16713, -32'd1421, -32'd8345, 32'd389},
{-32'd4769, -32'd1154, 32'd3648, -32'd1561},
{-32'd4844, 32'd178, 32'd11044, -32'd4242},
{-32'd3981, -32'd1160, 32'd4087, -32'd624},
{32'd15050, -32'd4243, 32'd9293, 32'd3242},
{-32'd18045, -32'd12789, 32'd9976, 32'd9824},
{32'd1200, 32'd9599, 32'd9569, 32'd5454},
{32'd957, 32'd6984, -32'd1586, -32'd6285},
{-32'd3403, 32'd2266, 32'd4259, 32'd4267},
{-32'd4005, -32'd2209, -32'd18801, -32'd5731},
{32'd3318, 32'd6438, -32'd4063, 32'd5317},
{-32'd5514, -32'd1203, -32'd2213, 32'd2724},
{-32'd8214, 32'd10042, 32'd3447, 32'd9309},
{32'd3751, 32'd7960, -32'd7001, 32'd3496},
{-32'd13084, 32'd522, 32'd1361, 32'd11602},
{-32'd2236, -32'd3936, 32'd8762, 32'd575},
{-32'd8877, 32'd13321, 32'd215, 32'd693},
{32'd4063, 32'd6863, 32'd7864, -32'd11279},
{-32'd1439, -32'd648, -32'd11432, -32'd7557},
{32'd6079, 32'd1905, -32'd10858, -32'd1911},
{-32'd789, 32'd324, 32'd7038, 32'd2465},
{32'd5837, -32'd1873, 32'd1175, 32'd9596},
{-32'd3423, 32'd2834, -32'd5492, -32'd8537},
{32'd6390, -32'd3149, 32'd7283, -32'd938},
{-32'd7497, 32'd5780, 32'd3306, 32'd11112},
{32'd2755, -32'd2006, 32'd632, 32'd4401},
{-32'd4760, 32'd9735, 32'd6896, 32'd7793},
{-32'd971, 32'd2579, -32'd3350, 32'd3395},
{-32'd11218, 32'd5549, 32'd7766, -32'd9848},
{-32'd2521, 32'd9705, -32'd1276, 32'd1464},
{-32'd16238, -32'd5268, -32'd1545, -32'd5448},
{32'd11963, -32'd1037, 32'd1013, 32'd4148},
{32'd2402, 32'd6530, -32'd421, -32'd11674},
{-32'd9944, 32'd252, -32'd5953, -32'd585},
{32'd7306, 32'd854, 32'd5832, -32'd3765},
{32'd1451, -32'd1476, -32'd1900, 32'd2867},
{32'd5874, 32'd4073, 32'd3632, 32'd1553},
{32'd6212, -32'd7595, -32'd1123, -32'd1371},
{-32'd16954, -32'd2806, 32'd4275, 32'd3921},
{32'd9111, -32'd2866, 32'd6573, -32'd4980},
{32'd1841, 32'd11632, 32'd18519, 32'd5948},
{-32'd11448, -32'd14471, 32'd84, 32'd3641},
{-32'd286, -32'd5972, -32'd3672, -32'd9863},
{-32'd2780, -32'd7299, 32'd16468, 32'd9620},
{-32'd8009, -32'd5058, 32'd3421, 32'd1685},
{-32'd2738, -32'd8144, -32'd9858, 32'd5558},
{-32'd8021, -32'd3682, 32'd9503, 32'd12576},
{32'd6358, 32'd5962, 32'd1845, 32'd4631},
{-32'd13130, 32'd1901, -32'd3359, -32'd7663},
{-32'd2410, -32'd12788, -32'd227, 32'd6666},
{-32'd1552, 32'd9051, 32'd3526, -32'd2956},
{-32'd5753, -32'd4082, -32'd1854, -32'd5732},
{32'd1174, -32'd1672, 32'd596, -32'd10323},
{32'd6998, 32'd3471, -32'd4566, -32'd3671},
{-32'd2505, -32'd7184, 32'd8523, -32'd3079},
{32'd3442, 32'd9649, 32'd5986, 32'd1732},
{32'd489, 32'd3739, -32'd13135, 32'd6228},
{32'd2877, 32'd5752, 32'd24, -32'd9539},
{32'd2158, 32'd5284, -32'd2756, -32'd11033},
{-32'd4102, -32'd2012, -32'd4214, 32'd4256},
{-32'd6336, 32'd231, -32'd5550, 32'd8287},
{32'd1234, 32'd2144, 32'd5562, 32'd577},
{32'd3124, 32'd13593, 32'd8823, 32'd4658},
{32'd1599, 32'd9181, -32'd11469, -32'd2643},
{-32'd7222, -32'd428, 32'd5102, -32'd7794},
{32'd2573, -32'd3433, 32'd40, 32'd5035},
{-32'd3865, 32'd4082, 32'd1355, -32'd870},
{32'd12267, 32'd2385, 32'd6967, -32'd654},
{-32'd3714, 32'd795, 32'd1382, -32'd3724},
{32'd1386, 32'd4413, -32'd7013, 32'd636},
{32'd4056, 32'd7231, 32'd1722, -32'd3097},
{-32'd6720, 32'd916, 32'd4970, 32'd6516},
{32'd1570, 32'd2500, -32'd7667, 32'd6394},
{32'd2013, 32'd449, 32'd14437, 32'd5585},
{-32'd381, 32'd3014, 32'd1394, 32'd6574},
{-32'd2248, -32'd477, 32'd17268, -32'd1568},
{-32'd14888, -32'd6000, -32'd6258, 32'd2930},
{32'd9802, -32'd5941, 32'd9536, 32'd6307},
{32'd9312, -32'd5005, 32'd4425, 32'd11261},
{32'd12314, 32'd1975, -32'd1722, 32'd538},
{-32'd2936, 32'd1375, -32'd8398, -32'd8113},
{-32'd7084, 32'd15219, 32'd5218, -32'd7984},
{32'd7383, -32'd10125, 32'd3155, 32'd4521},
{32'd5365, -32'd5799, 32'd12220, -32'd1055},
{32'd5349, 32'd366, 32'd7389, 32'd928},
{-32'd2457, 32'd11072, -32'd2119, -32'd5253},
{-32'd5197, 32'd627, -32'd4848, -32'd7217},
{32'd4140, -32'd4574, -32'd5421, 32'd6602},
{-32'd7244, -32'd2259, -32'd435, -32'd2346},
{-32'd11591, -32'd5835, 32'd5217, 32'd6036},
{-32'd2177, -32'd3097, 32'd8472, 32'd11261},
{32'd3432, -32'd10358, -32'd16431, -32'd1955},
{32'd422, 32'd1813, 32'd7416, -32'd4634},
{-32'd1126, -32'd3176, -32'd2774, 32'd2676},
{32'd10179, 32'd6919, 32'd12268, 32'd5416},
{32'd3342, 32'd1544, 32'd5066, -32'd921},
{-32'd10869, -32'd10028, -32'd12832, 32'd3506},
{-32'd716, 32'd9841, -32'd2615, -32'd6321},
{32'd9081, 32'd1787, 32'd5413, -32'd2205},
{32'd13453, 32'd4121, -32'd87, -32'd3909},
{32'd8596, 32'd3426, 32'd11295, 32'd4340},
{32'd4452, 32'd3854, -32'd13245, -32'd363},
{32'd4304, -32'd4541, -32'd1090, -32'd6508},
{-32'd7695, -32'd3485, -32'd3565, -32'd1756},
{32'd2243, -32'd4749, 32'd1563, 32'd2317},
{32'd3014, 32'd3217, -32'd4012, -32'd4781},
{32'd12838, 32'd3306, -32'd12565, -32'd636},
{32'd12277, -32'd2853, -32'd17993, -32'd810},
{-32'd11353, -32'd9570, 32'd7206, 32'd6053},
{32'd12328, 32'd4925, 32'd9312, -32'd458},
{-32'd891, 32'd1885, 32'd3863, 32'd3114},
{-32'd377, -32'd2404, -32'd10201, -32'd5989},
{-32'd1552, -32'd3276, -32'd5485, -32'd13527},
{-32'd7647, -32'd2590, -32'd4723, -32'd7183},
{32'd1211, 32'd10155, -32'd6013, 32'd6773},
{32'd4335, 32'd2852, 32'd699, -32'd3252},
{32'd4340, -32'd3893, 32'd5192, -32'd1322},
{-32'd7609, -32'd676, -32'd13546, -32'd1645}
},
{{32'd1737, 32'd7924, 32'd2639, 32'd5486},
{-32'd12603, -32'd2873, 32'd1490, -32'd7144},
{-32'd7528, -32'd4837, -32'd514, 32'd1281},
{32'd318, 32'd3896, 32'd5325, 32'd985},
{32'd335, -32'd5484, 32'd3721, -32'd3911},
{-32'd8633, 32'd6689, 32'd1484, 32'd1471},
{32'd795, -32'd562, 32'd413, -32'd3311},
{32'd6075, -32'd3392, 32'd8281, -32'd7272},
{-32'd132, 32'd3484, -32'd1325, 32'd3701},
{32'd9461, 32'd9550, 32'd4428, 32'd11616},
{-32'd5705, -32'd1653, 32'd695, 32'd2043},
{32'd9497, 32'd5029, 32'd2738, -32'd4478},
{32'd3046, 32'd2578, -32'd12779, 32'd9826},
{-32'd6808, 32'd1297, 32'd80, 32'd251},
{-32'd10212, -32'd10503, -32'd2064, 32'd2258},
{32'd13013, -32'd1268, -32'd7474, -32'd10869},
{32'd12022, 32'd114, 32'd19611, -32'd4502},
{32'd5116, 32'd837, -32'd2181, -32'd590},
{-32'd5522, -32'd290, -32'd3803, -32'd2353},
{32'd12057, 32'd9691, 32'd4942, 32'd1999},
{32'd3082, 32'd2132, -32'd10076, -32'd8035},
{-32'd16266, -32'd2260, -32'd2473, -32'd4345},
{-32'd1649, -32'd10511, -32'd4407, -32'd6136},
{-32'd6853, -32'd5134, -32'd5618, -32'd5454},
{32'd3387, 32'd8756, 32'd5321, 32'd5989},
{32'd3515, 32'd8405, -32'd3131, -32'd1432},
{32'd760, 32'd2578, 32'd298, 32'd10},
{-32'd4076, -32'd553, -32'd3723, -32'd228},
{32'd5125, -32'd6424, 32'd6916, -32'd4255},
{-32'd10177, 32'd447, -32'd5938, 32'd2388},
{-32'd1954, 32'd3116, 32'd3586, 32'd857},
{-32'd14607, 32'd5301, 32'd2298, -32'd3730},
{32'd8399, 32'd3597, 32'd7240, -32'd1691},
{-32'd6275, -32'd9390, -32'd6052, 32'd1377},
{32'd13321, 32'd6831, -32'd3203, 32'd4684},
{-32'd8347, 32'd3743, 32'd4049, -32'd565},
{32'd11635, 32'd6945, -32'd5387, 32'd520},
{32'd10304, -32'd3494, -32'd7335, -32'd3205},
{32'd2095, -32'd1535, 32'd10520, -32'd5026},
{-32'd2817, 32'd4055, -32'd316, -32'd717},
{32'd9284, 32'd3529, -32'd6051, 32'd2065},
{32'd9204, 32'd10941, 32'd2721, 32'd2773},
{32'd7050, 32'd2742, 32'd12102, 32'd1711},
{-32'd1841, -32'd12191, -32'd4604, -32'd4389},
{-32'd9730, -32'd2964, -32'd2199, -32'd3367},
{-32'd7195, 32'd2881, 32'd894, 32'd2623},
{-32'd3165, 32'd7062, -32'd8488, -32'd762},
{-32'd596, -32'd1105, 32'd3203, -32'd6303},
{32'd14485, 32'd3382, 32'd498, 32'd3673},
{-32'd2359, -32'd9641, -32'd2378, -32'd5819},
{32'd793, 32'd8889, 32'd8018, 32'd4034},
{32'd1662, 32'd1482, -32'd6336, 32'd775},
{-32'd6693, -32'd7208, 32'd3574, -32'd3258},
{32'd7014, 32'd98, -32'd2428, -32'd1301},
{32'd5457, -32'd297, -32'd1814, -32'd5334},
{-32'd2519, 32'd3153, 32'd3228, 32'd1719},
{32'd7250, 32'd8527, 32'd5276, -32'd2674},
{32'd2831, -32'd15236, -32'd1236, -32'd9138},
{32'd6563, -32'd12790, -32'd5636, -32'd1819},
{-32'd6472, 32'd5702, 32'd3337, -32'd5577},
{-32'd362, -32'd2635, 32'd4255, -32'd8447},
{-32'd2403, 32'd10775, -32'd3935, -32'd2481},
{-32'd2671, -32'd4912, 32'd2410, -32'd1152},
{-32'd3785, 32'd230, 32'd348, -32'd1562},
{-32'd2499, -32'd8380, -32'd3420, -32'd4738},
{-32'd3054, 32'd7338, 32'd4437, 32'd3984},
{32'd50, -32'd7675, -32'd1658, 32'd4789},
{-32'd6963, 32'd4001, -32'd6075, 32'd809},
{-32'd3241, -32'd11790, 32'd962, -32'd2931},
{32'd2655, -32'd2471, 32'd2177, -32'd3183},
{32'd999, -32'd5361, -32'd6466, -32'd1108},
{-32'd779, -32'd1575, -32'd5948, -32'd252},
{-32'd12156, 32'd2887, -32'd5874, -32'd2463},
{32'd1145, -32'd4492, 32'd1428, 32'd212},
{-32'd4765, -32'd1920, -32'd629, 32'd217},
{-32'd3058, -32'd4101, -32'd1932, -32'd2669},
{32'd801, -32'd12210, -32'd8463, -32'd5318},
{-32'd1256, -32'd10688, 32'd7992, -32'd2138},
{32'd4083, 32'd4929, 32'd380, 32'd7825},
{-32'd3062, -32'd3264, 32'd11436, 32'd532},
{32'd14747, 32'd10351, -32'd5245, -32'd6082},
{-32'd3058, -32'd6316, 32'd10003, 32'd2601},
{32'd4315, -32'd13721, 32'd1826, -32'd9820},
{32'd5267, -32'd477, -32'd3971, -32'd4433},
{-32'd2733, -32'd11373, 32'd5021, -32'd818},
{-32'd12179, 32'd5916, 32'd6841, -32'd1558},
{32'd5250, 32'd2921, -32'd634, 32'd6195},
{-32'd2748, -32'd12472, -32'd1747, -32'd7966},
{32'd8000, -32'd12405, 32'd11883, -32'd2618},
{32'd6147, -32'd3436, 32'd8489, -32'd3576},
{-32'd2388, 32'd5030, -32'd3127, 32'd742},
{-32'd1714, -32'd4464, 32'd1297, -32'd881},
{-32'd7273, 32'd4419, -32'd7915, 32'd8629},
{32'd5248, 32'd8962, -32'd8383, 32'd1771},
{32'd2521, -32'd8893, 32'd3361, -32'd3053},
{-32'd3476, -32'd2952, 32'd4129, 32'd1619},
{32'd1203, 32'd2760, -32'd1124, -32'd506},
{32'd8396, 32'd1648, 32'd2149, -32'd4751},
{32'd10340, -32'd364, 32'd3118, -32'd2058},
{32'd5194, 32'd6671, 32'd3181, 32'd1021},
{-32'd2281, -32'd12930, -32'd15009, -32'd1182},
{-32'd12896, -32'd2161, -32'd3016, -32'd2724},
{32'd1308, -32'd5926, -32'd4807, 32'd3553},
{32'd5830, -32'd9987, -32'd3735, 32'd3495},
{32'd6150, -32'd1550, -32'd309, 32'd3946},
{-32'd14989, 32'd5705, -32'd1049, -32'd2215},
{-32'd4983, 32'd2241, -32'd141, 32'd4045},
{-32'd5276, 32'd67, 32'd5261, 32'd1927},
{32'd4945, -32'd5459, 32'd1996, 32'd3554},
{32'd5809, 32'd3879, 32'd5265, -32'd7067},
{32'd4127, -32'd6027, -32'd3521, 32'd123},
{32'd11254, -32'd11784, 32'd5561, -32'd4641},
{32'd4219, 32'd1273, 32'd8264, 32'd5556},
{-32'd77, -32'd5130, 32'd4272, 32'd66},
{-32'd1198, -32'd482, 32'd4106, -32'd3082},
{32'd8187, -32'd4073, 32'd118, 32'd3683},
{-32'd7997, -32'd886, -32'd372, 32'd1056},
{-32'd6871, 32'd4637, -32'd8642, -32'd8497},
{32'd7526, 32'd2167, -32'd2794, -32'd7891},
{32'd647, 32'd14041, 32'd5027, 32'd12105},
{-32'd8290, 32'd554, 32'd2946, 32'd2152},
{-32'd3915, -32'd187, -32'd7934, -32'd2049},
{-32'd11660, 32'd2832, 32'd86, 32'd1997},
{-32'd11119, 32'd89, -32'd2005, -32'd2252},
{32'd5779, -32'd4498, 32'd3532, -32'd4063},
{-32'd5381, 32'd17324, 32'd8011, 32'd3761},
{-32'd4391, 32'd2061, 32'd8040, 32'd7984},
{-32'd9992, -32'd3066, -32'd12479, -32'd4691},
{32'd6223, -32'd2801, -32'd2805, -32'd3622},
{32'd7920, -32'd4288, -32'd622, -32'd5936},
{-32'd10667, 32'd3021, 32'd14295, 32'd2267},
{-32'd8258, -32'd8031, 32'd3754, -32'd2129},
{-32'd4262, -32'd2720, -32'd9958, -32'd232},
{-32'd10486, 32'd2160, -32'd6236, -32'd2454},
{-32'd7564, -32'd2826, -32'd465, -32'd3649},
{-32'd857, -32'd2087, 32'd2685, -32'd3208},
{-32'd3513, 32'd3922, -32'd11507, -32'd1137},
{-32'd6033, 32'd5765, -32'd3559, 32'd1266},
{32'd2681, -32'd7500, 32'd3861, -32'd1108},
{-32'd3651, -32'd9044, -32'd6107, -32'd7256},
{-32'd1069, -32'd957, 32'd9826, -32'd2153},
{32'd225, -32'd1229, -32'd2480, 32'd2307},
{-32'd15076, 32'd7371, 32'd1818, -32'd4931},
{32'd4369, 32'd6057, -32'd7398, -32'd2272},
{-32'd2652, 32'd3394, -32'd3466, 32'd5147},
{32'd14268, -32'd5743, 32'd12598, -32'd3533},
{-32'd430, -32'd5825, -32'd1213, -32'd1430},
{-32'd8629, -32'd1282, -32'd9407, 32'd8337},
{-32'd2524, 32'd3111, 32'd5537, 32'd252},
{-32'd11650, -32'd7776, 32'd8275, -32'd1692},
{32'd13, 32'd1941, -32'd9944, -32'd2887},
{32'd3432, 32'd9169, 32'd6820, 32'd1078},
{32'd15047, -32'd1098, 32'd4317, -32'd2172},
{32'd1123, 32'd3247, 32'd396, -32'd3701},
{32'd4468, -32'd5783, -32'd9751, -32'd253},
{-32'd2057, -32'd12057, -32'd6271, -32'd10162},
{32'd15005, 32'd3365, 32'd453, 32'd2757},
{-32'd872, 32'd5879, -32'd2558, -32'd1300},
{32'd10094, -32'd3423, -32'd8767, -32'd2889},
{32'd972, 32'd747, -32'd1749, 32'd7300},
{-32'd4226, -32'd6152, -32'd3881, -32'd4548},
{-32'd1007, -32'd4725, -32'd3441, -32'd772},
{-32'd749, -32'd4251, -32'd8261, -32'd5119},
{32'd266, 32'd1811, -32'd3892, 32'd284},
{32'd2900, 32'd3834, -32'd2062, -32'd1120},
{-32'd3366, -32'd7637, 32'd1339, 32'd5580},
{-32'd5540, 32'd3284, -32'd10678, 32'd7798},
{-32'd3879, -32'd4696, 32'd5757, -32'd5786},
{32'd199, -32'd1584, 32'd986, 32'd386},
{-32'd449, -32'd6028, 32'd7359, -32'd941},
{-32'd346, -32'd120, -32'd9521, 32'd4694},
{32'd941, -32'd3840, -32'd3423, -32'd1095},
{32'd8204, 32'd5318, 32'd5443, 32'd4746},
{-32'd9213, -32'd180, -32'd5383, -32'd525},
{-32'd3857, 32'd6076, -32'd5364, 32'd2484},
{32'd12779, -32'd841, -32'd193, 32'd7967},
{32'd757, 32'd6892, 32'd13504, -32'd3745},
{-32'd5618, 32'd2173, -32'd9375, 32'd4253},
{-32'd772, 32'd1103, -32'd212, -32'd2869},
{-32'd4715, 32'd247, 32'd4179, -32'd5924},
{32'd2278, -32'd6373, -32'd7254, -32'd2336},
{-32'd3823, -32'd1673, 32'd1110, 32'd395},
{-32'd5851, -32'd6100, 32'd3370, 32'd1834},
{-32'd3376, -32'd6957, 32'd425, 32'd1997},
{32'd2137, -32'd6760, -32'd3318, 32'd1966},
{32'd12092, 32'd14098, 32'd7391, 32'd6101},
{32'd2225, 32'd7361, -32'd4071, 32'd1946},
{-32'd4506, -32'd61, 32'd1157, 32'd623},
{-32'd131, -32'd1455, -32'd8694, -32'd3829},
{-32'd219, -32'd761, 32'd2556, -32'd7078},
{32'd1107, 32'd5180, -32'd9717, -32'd2146},
{-32'd4951, -32'd59, 32'd2796, 32'd2682},
{32'd3189, -32'd13, 32'd579, -32'd837},
{-32'd5567, 32'd5175, -32'd10877, 32'd7385},
{-32'd6198, -32'd2861, 32'd4863, 32'd6607},
{32'd2758, -32'd2237, 32'd379, -32'd4677},
{32'd504, -32'd11397, -32'd7755, -32'd2356},
{-32'd2629, 32'd4360, 32'd3541, 32'd5936},
{32'd2235, 32'd13020, -32'd7900, -32'd4482},
{32'd8026, -32'd1143, -32'd5475, -32'd3372},
{-32'd4075, -32'd4511, -32'd6325, -32'd3480},
{-32'd4012, -32'd2894, 32'd220, -32'd80},
{-32'd1448, -32'd391, -32'd31, -32'd6434},
{32'd9337, 32'd10638, 32'd4078, 32'd2665},
{32'd2822, -32'd14944, -32'd8907, -32'd4592},
{32'd4178, 32'd2288, -32'd5882, -32'd936},
{-32'd8149, -32'd802, -32'd1070, 32'd12537},
{-32'd3278, -32'd11878, 32'd5884, -32'd7391},
{32'd14046, -32'd4195, -32'd537, 32'd4386},
{-32'd6400, -32'd4637, -32'd1387, -32'd2264},
{32'd7790, -32'd2771, -32'd12945, 32'd6222},
{-32'd1772, -32'd3301, -32'd9262, 32'd5777},
{-32'd4633, 32'd2909, 32'd2688, -32'd2771},
{32'd9155, -32'd1367, -32'd3239, 32'd9095},
{-32'd3542, 32'd680, -32'd3610, -32'd1331},
{-32'd9261, 32'd7414, -32'd106, -32'd2267},
{32'd3679, 32'd943, 32'd1878, -32'd8744},
{-32'd5861, -32'd95, 32'd1508, -32'd1446},
{-32'd175, -32'd730, -32'd1800, -32'd1689},
{-32'd10462, -32'd7040, -32'd3799, -32'd5256},
{32'd3206, -32'd5947, -32'd783, 32'd502},
{-32'd356, -32'd5596, 32'd7522, -32'd1576},
{32'd5873, -32'd1155, -32'd1586, -32'd1329},
{-32'd670, -32'd1882, -32'd5149, 32'd2208},
{32'd815, 32'd7338, 32'd1733, -32'd4529},
{-32'd1271, 32'd1688, -32'd19, -32'd5211},
{32'd1664, -32'd4263, -32'd1581, -32'd303},
{-32'd7418, 32'd6245, 32'd13594, -32'd6367},
{32'd8723, -32'd2091, 32'd6015, 32'd639},
{-32'd8243, -32'd1589, 32'd7354, 32'd2486},
{32'd5092, -32'd1459, -32'd9619, -32'd2431},
{-32'd8201, 32'd477, 32'd4705, -32'd6074},
{32'd7656, 32'd9893, -32'd1595, 32'd4187},
{-32'd4696, -32'd3737, -32'd8560, 32'd947},
{-32'd4102, 32'd30, -32'd3003, 32'd2324},
{-32'd8320, -32'd14512, 32'd65, 32'd621},
{32'd1665, -32'd8014, 32'd2082, 32'd3318},
{-32'd3270, 32'd6844, 32'd252, 32'd3380},
{32'd3270, -32'd325, 32'd11425, -32'd1292},
{-32'd4257, -32'd5242, 32'd2337, -32'd8955},
{-32'd451, 32'd4274, -32'd1050, -32'd4937},
{32'd845, -32'd2682, 32'd473, 32'd3174},
{-32'd11492, -32'd3771, -32'd9413, -32'd5201},
{-32'd6207, 32'd2732, -32'd621, 32'd4003},
{32'd16626, 32'd6536, 32'd4475, 32'd4915},
{32'd459, -32'd3047, -32'd2981, -32'd4258},
{32'd6252, -32'd100, 32'd132, -32'd5091},
{-32'd4833, 32'd7230, 32'd11524, 32'd556},
{32'd7268, -32'd2361, 32'd425, 32'd748},
{-32'd13998, -32'd2213, -32'd1536, 32'd1124},
{32'd1195, -32'd11583, 32'd12147, -32'd2032},
{-32'd2288, -32'd6690, 32'd4469, 32'd4759},
{32'd1281, -32'd598, 32'd106, -32'd4675},
{-32'd1839, 32'd9356, -32'd1122, -32'd305},
{32'd2732, -32'd6344, -32'd7675, -32'd1309},
{32'd8082, 32'd4479, -32'd1080, -32'd1127},
{32'd5043, 32'd5594, 32'd2523, -32'd614},
{-32'd2217, 32'd9736, 32'd7882, 32'd2808},
{32'd1030, -32'd18641, -32'd2546, -32'd1871},
{32'd1349, 32'd3645, 32'd2608, -32'd267},
{32'd5820, 32'd8324, -32'd1537, -32'd1331},
{32'd12088, 32'd749, 32'd3237, -32'd4294},
{-32'd7698, -32'd545, -32'd1697, -32'd37},
{-32'd1941, -32'd7697, -32'd1926, -32'd574},
{32'd7833, 32'd9415, -32'd12322, 32'd7006},
{-32'd2083, -32'd7601, 32'd7268, -32'd2893},
{32'd2261, 32'd12846, 32'd9379, 32'd83},
{32'd835, -32'd6231, -32'd7575, 32'd1899},
{32'd5859, -32'd17981, 32'd1892, -32'd1846},
{32'd12, -32'd3682, 32'd5963, -32'd7364},
{-32'd1991, -32'd12541, -32'd2893, -32'd38},
{32'd922, -32'd899, 32'd4860, 32'd4037},
{32'd8360, 32'd3989, 32'd1347, -32'd1740},
{-32'd2225, 32'd1122, -32'd7667, 32'd1940},
{-32'd11331, 32'd120, 32'd3387, -32'd1686},
{32'd11570, 32'd1068, -32'd7973, -32'd1759},
{32'd9622, 32'd8433, 32'd5839, 32'd5996},
{32'd4389, 32'd2310, -32'd186, 32'd2804},
{-32'd7484, -32'd4844, 32'd2938, -32'd10138},
{-32'd6928, 32'd7654, -32'd4015, -32'd781},
{-32'd1033, 32'd846, -32'd7657, 32'd3976},
{32'd3539, 32'd2918, 32'd4738, 32'd2160},
{32'd14412, 32'd3957, -32'd1126, -32'd4606},
{-32'd11491, 32'd6146, 32'd3355, 32'd3157},
{32'd10977, 32'd10100, -32'd1324, -32'd4897},
{-32'd7541, -32'd8214, -32'd1277, -32'd8407},
{32'd1198, -32'd1944, 32'd6867, 32'd2815},
{32'd5186, 32'd3922, -32'd2333, 32'd6308},
{-32'd1029, 32'd776, -32'd6624, -32'd3149},
{-32'd2374, 32'd8127, 32'd7595, -32'd2086},
{-32'd851, 32'd56, -32'd7222, 32'd1609},
{32'd4283, 32'd14254, 32'd1177, 32'd2827},
{32'd6711, 32'd5369, 32'd5184, -32'd4837},
{-32'd9194, -32'd2570, -32'd4740, 32'd365},
{-32'd8130, -32'd2297, -32'd4312, 32'd164},
{32'd8257, -32'd1998, 32'd582, -32'd1926},
{-32'd3183, 32'd3480, 32'd178, -32'd2659},
{-32'd961, -32'd2392, 32'd3562, 32'd6887},
{-32'd2582, 32'd8210, 32'd7118, 32'd7592},
{32'd5593, -32'd12362, 32'd814, -32'd7882}
},
{{32'd5017, -32'd1343, -32'd28, 32'd3680},
{32'd6057, -32'd27871, -32'd16672, -32'd17487},
{-32'd7235, -32'd1886, -32'd2618, 32'd7199},
{-32'd927, -32'd657, 32'd10109, 32'd5036},
{32'd4973, 32'd11599, -32'd8816, -32'd8610},
{32'd2562, -32'd6881, 32'd2588, 32'd1489},
{32'd5303, 32'd12373, 32'd4554, 32'd12448},
{32'd3878, -32'd3527, 32'd13885, -32'd6528},
{32'd16097, -32'd3765, 32'd975, 32'd1461},
{32'd5019, -32'd493, 32'd10628, 32'd8166},
{-32'd6080, -32'd12253, -32'd3381, -32'd925},
{32'd5342, 32'd1393, -32'd2389, -32'd8075},
{32'd18559, -32'd530, -32'd11840, -32'd808},
{32'd3412, 32'd248, -32'd8942, -32'd11756},
{-32'd2918, 32'd1767, 32'd4587, -32'd4617},
{32'd1941, -32'd3355, -32'd8236, -32'd883},
{32'd18908, 32'd5786, 32'd1066, 32'd5027},
{-32'd23311, -32'd12585, 32'd2646, -32'd7556},
{32'd2812, 32'd9671, 32'd4015, -32'd2940},
{32'd27417, -32'd9188, -32'd4404, 32'd8870},
{32'd14744, 32'd3401, 32'd4422, 32'd4604},
{-32'd1130, 32'd3847, 32'd3414, -32'd2653},
{32'd8390, -32'd8320, 32'd343, -32'd11454},
{-32'd19914, 32'd3198, 32'd12360, -32'd1048},
{-32'd6156, -32'd4001, 32'd7111, 32'd355},
{-32'd16649, 32'd18483, -32'd6978, -32'd4961},
{-32'd8684, -32'd1440, 32'd4871, -32'd323},
{-32'd3035, -32'd2832, 32'd3290, -32'd1795},
{32'd4001, -32'd14482, -32'd9582, -32'd7857},
{-32'd16156, 32'd8317, -32'd4181, 32'd10357},
{32'd4628, -32'd1791, 32'd4117, -32'd10504},
{-32'd6408, -32'd4805, -32'd5058, -32'd15510},
{32'd8210, 32'd13169, 32'd2780, -32'd1606},
{-32'd19838, 32'd8969, -32'd12007, -32'd6746},
{32'd4642, 32'd5958, 32'd12226, 32'd15086},
{32'd7371, 32'd8631, 32'd2049, 32'd2818},
{-32'd7178, -32'd669, 32'd10086, 32'd4187},
{32'd2944, -32'd1776, -32'd5931, -32'd7853},
{-32'd5521, -32'd11713, -32'd654, 32'd7686},
{-32'd12910, 32'd4433, 32'd2348, 32'd1943},
{-32'd6094, -32'd34, -32'd21000, -32'd1817},
{-32'd916, 32'd4397, 32'd836, -32'd2387},
{-32'd6383, 32'd3231, -32'd2795, -32'd736},
{32'd4932, 32'd10156, -32'd15006, -32'd8668},
{-32'd1436, 32'd10443, 32'd9, 32'd2248},
{-32'd472, -32'd4482, -32'd15886, 32'd47},
{-32'd59, -32'd3875, 32'd8274, -32'd7747},
{-32'd10226, 32'd8896, -32'd10989, -32'd940},
{32'd6839, -32'd7648, 32'd3213, 32'd6885},
{32'd4331, 32'd376, 32'd562, -32'd12088},
{-32'd2669, -32'd9210, 32'd2698, -32'd2290},
{-32'd11247, -32'd3385, -32'd2416, -32'd9661},
{-32'd2261, 32'd6728, 32'd2034, 32'd897},
{32'd5894, 32'd15243, 32'd1426, -32'd492},
{-32'd1704, 32'd5407, -32'd7792, 32'd1486},
{32'd3346, -32'd12464, 32'd2335, -32'd9964},
{-32'd8981, 32'd4184, -32'd924, 32'd8783},
{-32'd17773, 32'd1381, -32'd2526, -32'd3273},
{-32'd5898, 32'd2072, -32'd480, -32'd10504},
{-32'd1398, -32'd3604, 32'd3328, 32'd784},
{32'd11235, 32'd10606, -32'd2249, -32'd4130},
{-32'd6724, 32'd3169, 32'd2231, 32'd6854},
{32'd5002, -32'd13879, -32'd4131, -32'd7993},
{32'd8525, 32'd1758, -32'd7006, -32'd6680},
{-32'd9679, -32'd11611, -32'd13605, 32'd6376},
{32'd6037, 32'd2447, 32'd19444, 32'd12761},
{32'd3457, 32'd7125, -32'd11134, -32'd3128},
{-32'd1936, -32'd25120, -32'd5914, -32'd4450},
{-32'd429, -32'd5109, -32'd1320, -32'd4534},
{-32'd2057, 32'd5631, 32'd750, 32'd7230},
{32'd1796, -32'd5678, -32'd3054, -32'd3427},
{32'd6243, 32'd7035, 32'd7973, -32'd10779},
{-32'd285, 32'd14393, -32'd2383, -32'd3677},
{32'd1266, 32'd3622, -32'd6653, 32'd6413},
{32'd4017, 32'd8673, 32'd37, 32'd722},
{-32'd20553, 32'd10360, 32'd89, -32'd292},
{-32'd5996, -32'd2992, -32'd6804, -32'd6149},
{-32'd15449, 32'd4688, -32'd2992, -32'd2191},
{32'd6144, 32'd11981, 32'd4310, 32'd6883},
{-32'd7739, 32'd3189, 32'd9786, 32'd10547},
{-32'd18833, -32'd4115, 32'd1321, -32'd3161},
{32'd10150, 32'd6328, 32'd8053, -32'd3680},
{32'd1573, 32'd4749, 32'd3205, 32'd3909},
{-32'd11019, -32'd3796, -32'd3993, -32'd9941},
{-32'd21158, 32'd4541, -32'd2945, -32'd5084},
{32'd4299, 32'd14857, -32'd12361, -32'd7015},
{-32'd2446, -32'd956, -32'd3939, 32'd3181},
{32'd2970, -32'd4199, 32'd11533, -32'd1065},
{32'd1816, -32'd2222, -32'd4557, 32'd4648},
{-32'd3051, 32'd10163, -32'd20217, -32'd2041},
{32'd1460, -32'd10255, -32'd7593, -32'd10688},
{-32'd513, -32'd6980, -32'd3874, 32'd30},
{32'd5164, 32'd1040, 32'd6896, -32'd1379},
{32'd176, -32'd12887, -32'd2041, -32'd1489},
{-32'd2006, 32'd13660, 32'd2149, -32'd7705},
{-32'd12513, -32'd19870, 32'd2494, -32'd9025},
{32'd3253, 32'd6006, 32'd14055, 32'd4916},
{-32'd6097, 32'd3502, 32'd6129, 32'd79},
{32'd2606, -32'd6078, 32'd3582, 32'd15472},
{-32'd1688, 32'd10496, 32'd12804, 32'd6777},
{32'd19170, -32'd3249, -32'd9790, -32'd8357},
{32'd1940, -32'd5866, -32'd3574, 32'd8491},
{-32'd8132, 32'd10616, -32'd6351, 32'd5803},
{32'd4401, 32'd4906, 32'd3339, 32'd11530},
{32'd7247, -32'd1956, 32'd2326, 32'd3612},
{-32'd7694, 32'd6593, 32'd7768, 32'd1673},
{32'd7661, -32'd5988, -32'd4246, -32'd7987},
{32'd8815, 32'd3063, -32'd8527, -32'd2781},
{32'd12393, -32'd8507, 32'd9483, 32'd5253},
{32'd2560, -32'd14798, -32'd8970, 32'd2410},
{-32'd17776, -32'd4934, 32'd10254, 32'd10481},
{-32'd695, 32'd3557, 32'd3750, 32'd6678},
{-32'd869, -32'd22, -32'd1410, 32'd8079},
{32'd2321, 32'd692, 32'd6974, 32'd2893},
{32'd9894, 32'd2723, -32'd8343, -32'd4787},
{32'd4819, -32'd14929, 32'd3385, -32'd6568},
{32'd7915, 32'd2810, 32'd1241, 32'd1995},
{32'd6327, -32'd8187, -32'd3541, -32'd4384},
{-32'd4482, -32'd5389, 32'd3639, -32'd559},
{32'd9294, -32'd3112, 32'd7302, -32'd2},
{32'd17642, 32'd12693, 32'd5772, -32'd1275},
{-32'd6756, 32'd14788, 32'd11214, -32'd13464},
{32'd9825, -32'd3656, -32'd3988, -32'd5050},
{32'd1955, 32'd490, 32'd8550, 32'd4435},
{-32'd2241, 32'd493, -32'd7271, 32'd5915},
{-32'd4885, -32'd13834, 32'd9857, -32'd2428},
{-32'd7931, 32'd1030, -32'd7040, -32'd9570},
{-32'd3221, -32'd8831, 32'd8083, -32'd924},
{32'd1395, -32'd7646, -32'd2925, 32'd1283},
{32'd4847, 32'd14815, 32'd9837, 32'd663},
{-32'd1419, 32'd860, 32'd989, 32'd705},
{32'd2494, -32'd3771, -32'd6676, -32'd2234},
{-32'd2123, 32'd7107, -32'd11439, 32'd6784},
{-32'd2336, -32'd8590, 32'd6304, -32'd1677},
{32'd7059, 32'd3336, 32'd9754, 32'd6701},
{32'd8522, 32'd5186, 32'd7515, -32'd3290},
{32'd11204, 32'd11148, -32'd1857, 32'd5407},
{-32'd8787, -32'd14085, -32'd1312, 32'd7217},
{32'd2793, 32'd1339, 32'd2227, -32'd2823},
{32'd3793, -32'd6910, -32'd16050, -32'd20758},
{32'd8239, -32'd1926, 32'd6443, -32'd885},
{-32'd5832, 32'd7422, 32'd3351, -32'd6013},
{-32'd11646, 32'd1506, -32'd1499, -32'd4051},
{32'd14443, -32'd11258, -32'd16620, -32'd8693},
{-32'd190, -32'd4051, 32'd6815, 32'd11354},
{32'd1398, -32'd13422, 32'd2360, -32'd2969},
{-32'd7026, -32'd14762, -32'd8536, -32'd5320},
{32'd7117, -32'd2266, 32'd8808, 32'd8596},
{32'd2813, 32'd90, 32'd15902, 32'd1551},
{-32'd153, 32'd1339, -32'd5106, -32'd11254},
{-32'd10203, -32'd1813, -32'd8760, -32'd8129},
{32'd8103, -32'd11889, 32'd5809, -32'd4030},
{32'd15388, -32'd2436, -32'd6061, -32'd2223},
{32'd10095, 32'd55, -32'd7393, -32'd5381},
{-32'd5127, 32'd2051, -32'd2134, -32'd1144},
{-32'd17936, 32'd10544, 32'd11953, 32'd4518},
{32'd7559, -32'd2596, -32'd1764, 32'd12492},
{-32'd4062, 32'd10016, 32'd1782, 32'd16565},
{-32'd7143, -32'd10485, -32'd4951, -32'd190},
{32'd24853, 32'd10797, -32'd1692, -32'd5309},
{32'd7108, 32'd509, 32'd5563, -32'd11303},
{32'd3287, 32'd3878, 32'd6346, -32'd2261},
{32'd9220, -32'd6616, 32'd955, -32'd7535},
{32'd7837, 32'd16785, 32'd9665, 32'd967},
{32'd363, -32'd8104, -32'd16679, 32'd12686},
{-32'd5618, -32'd5301, -32'd8556, -32'd606},
{-32'd189, 32'd620, 32'd1771, 32'd5651},
{-32'd7917, 32'd2838, -32'd1427, -32'd1517},
{-32'd11211, -32'd779, -32'd11049, 32'd3602},
{-32'd587, -32'd8324, -32'd13165, -32'd5797},
{-32'd9291, 32'd2671, -32'd6697, -32'd5549},
{32'd1850, -32'd304, 32'd534, 32'd3268},
{32'd997, 32'd4229, 32'd6373, 32'd15011},
{-32'd14344, 32'd1066, 32'd8833, -32'd99},
{32'd3652, 32'd3424, 32'd16978, -32'd4235},
{32'd9312, 32'd248, -32'd941, -32'd1577},
{32'd5953, 32'd10976, -32'd3330, 32'd465},
{32'd5514, -32'd3052, 32'd1122, 32'd1737},
{32'd13896, 32'd6810, 32'd7797, 32'd1054},
{-32'd11915, 32'd2210, -32'd2038, -32'd9177},
{-32'd14533, -32'd6132, -32'd8907, -32'd9178},
{32'd6806, 32'd6436, -32'd13802, -32'd5080},
{-32'd6241, -32'd7681, 32'd590, -32'd10268},
{32'd8064, -32'd10462, -32'd7895, -32'd13829},
{-32'd4620, 32'd4820, 32'd4967, 32'd2546},
{32'd10953, 32'd4948, -32'd790, -32'd1540},
{32'd8385, 32'd1722, 32'd8639, 32'd10261},
{32'd9368, -32'd12298, 32'd10733, -32'd5100},
{32'd10968, -32'd806, 32'd6385, 32'd3664},
{-32'd3315, 32'd17988, -32'd8781, -32'd3424},
{32'd8702, 32'd11511, -32'd4395, -32'd863},
{-32'd3960, 32'd5940, 32'd1804, -32'd7650},
{-32'd13556, -32'd6316, -32'd15859, 32'd655},
{32'd2151, -32'd4243, 32'd8449, 32'd11444},
{-32'd19403, -32'd11967, -32'd473, 32'd6311},
{-32'd13371, -32'd1658, -32'd883, 32'd1099},
{-32'd499, 32'd3184, -32'd6521, 32'd4578},
{32'd419, -32'd1855, 32'd3104, 32'd7551},
{-32'd7925, 32'd783, 32'd1023, -32'd4327},
{-32'd6070, -32'd7890, 32'd5696, -32'd9062},
{-32'd1811, -32'd5162, -32'd13668, -32'd12082},
{-32'd22231, 32'd5349, -32'd3278, 32'd6052},
{32'd15553, -32'd11261, 32'd6489, 32'd10987},
{32'd6913, -32'd7994, 32'd7450, -32'd1839},
{-32'd15973, -32'd1696, -32'd4472, -32'd9988},
{-32'd12298, -32'd14261, -32'd9007, 32'd5390},
{32'd19706, -32'd2817, 32'd9726, -32'd442},
{-32'd6384, -32'd5548, -32'd1792, -32'd9344},
{-32'd2518, 32'd500, 32'd5939, 32'd11734},
{-32'd14681, 32'd10630, -32'd5408, 32'd6529},
{-32'd2088, -32'd3560, -32'd13619, -32'd11786},
{-32'd314, -32'd16819, -32'd2194, 32'd2244},
{32'd7172, 32'd714, -32'd9165, -32'd8722},
{-32'd12863, -32'd4572, 32'd3121, -32'd1743},
{-32'd8300, -32'd3760, -32'd12619, -32'd5183},
{32'd658, -32'd10571, 32'd2394, -32'd6390},
{32'd12457, -32'd16132, 32'd8813, -32'd2758},
{-32'd9716, 32'd9427, -32'd5824, 32'd2751},
{32'd14109, -32'd3314, 32'd2162, 32'd12445},
{-32'd8857, 32'd13828, -32'd2940, -32'd5041},
{32'd7895, -32'd12473, 32'd3973, -32'd9053},
{32'd1430, 32'd8960, 32'd12189, -32'd5205},
{-32'd4423, 32'd7044, 32'd11874, -32'd6336},
{32'd12252, 32'd9512, -32'd681, 32'd2772},
{32'd2960, 32'd7826, -32'd8093, 32'd10880},
{32'd501, -32'd1507, -32'd4874, -32'd2358},
{32'd3986, -32'd110, -32'd3002, -32'd8078},
{-32'd5192, 32'd11543, 32'd14077, -32'd4481},
{-32'd1499, 32'd16368, 32'd7447, 32'd2253},
{32'd2032, -32'd7976, -32'd7, 32'd4641},
{-32'd7722, -32'd3137, -32'd6458, -32'd3854},
{32'd13929, 32'd3153, 32'd4795, -32'd2709},
{32'd2347, 32'd8053, -32'd1111, -32'd7459},
{-32'd469, 32'd8907, 32'd14020, -32'd1031},
{32'd1238, -32'd1490, 32'd949, -32'd13236},
{-32'd159, -32'd6839, 32'd3906, -32'd8191},
{32'd8102, -32'd14226, -32'd11708, 32'd9068},
{-32'd14986, 32'd4480, -32'd17860, -32'd3746},
{-32'd4547, 32'd3682, -32'd3586, 32'd12612},
{-32'd6940, 32'd10804, 32'd1683, -32'd3608},
{-32'd10053, 32'd13474, 32'd7850, 32'd10178},
{-32'd2201, 32'd2303, -32'd5841, -32'd3958},
{-32'd8408, 32'd6469, -32'd7167, -32'd8689},
{-32'd12313, -32'd706, 32'd5675, 32'd7469},
{32'd1535, -32'd4727, 32'd5033, 32'd9849},
{-32'd11596, 32'd10035, 32'd12811, 32'd762},
{-32'd11623, -32'd2296, -32'd549, -32'd11574},
{-32'd8404, -32'd2386, 32'd3303, -32'd6182},
{-32'd4263, 32'd5861, 32'd2189, -32'd10328},
{32'd9826, -32'd7009, -32'd8095, 32'd10313},
{32'd198, -32'd10035, -32'd4120, -32'd10229},
{32'd14432, 32'd6434, 32'd8020, -32'd906},
{-32'd10729, 32'd9109, 32'd4237, 32'd594},
{32'd21135, -32'd1779, 32'd9686, -32'd716},
{32'd233, -32'd8287, -32'd10110, -32'd10804},
{32'd8424, -32'd4199, 32'd3648, 32'd8515},
{32'd7872, -32'd7234, -32'd10060, 32'd325},
{-32'd6557, 32'd13495, 32'd14903, 32'd8484},
{32'd3833, 32'd11401, 32'd2499, -32'd6042},
{-32'd2431, -32'd12024, 32'd6090, 32'd2401},
{32'd2914, -32'd14613, 32'd4294, -32'd2672},
{-32'd9208, 32'd6333, -32'd9744, 32'd1099},
{-32'd18043, 32'd4720, -32'd5140, -32'd6812},
{-32'd9319, 32'd4484, 32'd3645, -32'd3872},
{32'd7429, -32'd5333, -32'd3127, 32'd2523},
{32'd11342, -32'd4012, -32'd8493, -32'd5467},
{32'd986, 32'd11117, 32'd5077, 32'd8625},
{-32'd8202, 32'd4117, 32'd2881, 32'd3477},
{-32'd2544, -32'd5705, -32'd4271, 32'd1151},
{32'd7528, -32'd11132, -32'd14275, 32'd1301},
{32'd881, -32'd10609, 32'd9549, 32'd5228},
{-32'd16643, -32'd1840, 32'd13270, 32'd6716},
{-32'd4898, -32'd8111, -32'd21535, -32'd10654},
{32'd8781, -32'd3078, -32'd164, -32'd6396},
{32'd9293, -32'd3853, 32'd4556, -32'd7974},
{32'd31, 32'd4869, -32'd6339, -32'd4177},
{32'd8526, 32'd2450, 32'd13133, 32'd8122},
{-32'd2791, -32'd18789, -32'd6111, 32'd10806},
{-32'd1078, 32'd10471, -32'd5776, -32'd10016},
{-32'd7246, 32'd6267, -32'd8435, 32'd3300},
{32'd14324, 32'd19508, 32'd7319, -32'd4621},
{32'd12812, -32'd19288, -32'd1691, -32'd9520},
{32'd2489, -32'd10059, -32'd7494, -32'd8528},
{32'd3019, -32'd8011, 32'd8656, 32'd4919},
{-32'd4972, -32'd1288, 32'd3512, 32'd4961},
{-32'd13871, -32'd7798, -32'd6839, -32'd5055},
{32'd3605, -32'd2884, 32'd10301, 32'd14729},
{-32'd14184, -32'd4926, -32'd3347, -32'd7742},
{32'd4155, -32'd699, 32'd13391, -32'd1706},
{-32'd1949, 32'd2376, 32'd3101, -32'd5972},
{32'd7381, -32'd4146, -32'd1409, 32'd4245},
{32'd3518, -32'd3459, 32'd16271, 32'd10192},
{-32'd5361, -32'd2153, -32'd5541, -32'd2471},
{-32'd4822, 32'd11894, -32'd11649, 32'd214},
{-32'd3829, -32'd1756, -32'd9064, -32'd5518},
{-32'd8083, 32'd1830, -32'd616, -32'd8294},
{-32'd2275, 32'd5707, -32'd5684, -32'd121},
{32'd4222, 32'd1083, 32'd8139, -32'd1011},
{-32'd6994, 32'd7662, 32'd13434, 32'd17642},
{32'd8085, 32'd1722, -32'd2321, -32'd705}
},
{{-32'd8411, 32'd2209, 32'd7185, -32'd179},
{-32'd18675, -32'd11643, -32'd13273, -32'd4714},
{-32'd2835, -32'd4816, -32'd2359, 32'd88},
{32'd14172, -32'd1206, -32'd1313, 32'd8138},
{-32'd128, 32'd4290, 32'd17266, 32'd2239},
{-32'd8758, 32'd5262, -32'd3538, 32'd4993},
{32'd8335, 32'd15577, 32'd10817, 32'd4231},
{32'd7882, 32'd1535, -32'd3055, -32'd5409},
{32'd12389, -32'd3557, 32'd16913, -32'd4482},
{32'd2134, 32'd10069, 32'd7358, -32'd17},
{-32'd6169, 32'd3225, -32'd3777, -32'd7636},
{-32'd4254, 32'd6387, 32'd204, -32'd2630},
{32'd8759, 32'd23388, 32'd5581, 32'd6244},
{-32'd11995, -32'd6184, -32'd6269, 32'd2299},
{32'd7815, 32'd6847, -32'd13276, -32'd4436},
{-32'd2525, -32'd3129, -32'd2755, -32'd5646},
{32'd1007, 32'd5231, -32'd3991, 32'd3515},
{-32'd3419, 32'd7560, 32'd4296, -32'd7766},
{-32'd2471, -32'd1320, 32'd5688, 32'd2543},
{-32'd4914, -32'd5950, 32'd4556, -32'd6631},
{32'd57, 32'd2397, 32'd10508, -32'd1657},
{-32'd9043, -32'd9994, -32'd5801, 32'd2715},
{-32'd3224, -32'd3505, -32'd1710, -32'd2392},
{-32'd824, 32'd2446, -32'd3281, 32'd3697},
{-32'd5993, 32'd8230, 32'd1738, -32'd6347},
{32'd1018, 32'd6355, 32'd598, 32'd4083},
{32'd6894, -32'd4979, 32'd9337, 32'd14827},
{32'd17539, 32'd15435, 32'd5727, -32'd4466},
{-32'd5969, 32'd11630, 32'd8393, 32'd2043},
{32'd3766, 32'd1300, 32'd1579, 32'd1469},
{-32'd5, 32'd3173, 32'd503, 32'd5552},
{-32'd6598, -32'd948, -32'd11551, -32'd545},
{32'd14493, 32'd3242, 32'd4940, -32'd6236},
{32'd10053, 32'd5047, -32'd1864, -32'd2996},
{32'd7022, 32'd10563, 32'd7299, 32'd1733},
{-32'd5875, -32'd9047, -32'd6049, 32'd4898},
{32'd4549, -32'd27, -32'd2260, -32'd4160},
{-32'd1156, -32'd15006, 32'd3698, -32'd2461},
{-32'd6373, -32'd437, 32'd4872, 32'd9287},
{32'd5318, 32'd6877, 32'd4878, -32'd1467},
{-32'd6972, -32'd4634, -32'd2157, -32'd714},
{32'd3533, 32'd9468, -32'd1707, 32'd5883},
{32'd2292, 32'd5576, 32'd3299, 32'd5772},
{-32'd2742, 32'd9708, 32'd1511, 32'd4623},
{32'd783, -32'd13427, 32'd5265, 32'd3893},
{32'd10424, -32'd1204, 32'd13813, 32'd3006},
{32'd121, 32'd2489, 32'd8184, 32'd2254},
{-32'd588, 32'd2772, 32'd88, 32'd3741},
{-32'd12087, 32'd9314, -32'd8579, 32'd91},
{-32'd18311, -32'd2710, -32'd174, -32'd5507},
{-32'd6152, -32'd13028, -32'd1076, -32'd6746},
{-32'd9595, 32'd5834, -32'd8094, 32'd953},
{-32'd3314, -32'd226, -32'd1650, -32'd5780},
{-32'd3606, 32'd9829, -32'd5978, 32'd430},
{32'd3669, 32'd15366, 32'd7109, 32'd1024},
{-32'd3657, -32'd1579, 32'd956, -32'd2396},
{-32'd13161, 32'd9084, 32'd7970, -32'd713},
{32'd7849, -32'd7665, -32'd16601, -32'd4404},
{32'd536, -32'd2472, -32'd11078, 32'd3994},
{32'd2845, 32'd10791, -32'd4495, -32'd6543},
{32'd6647, -32'd4802, 32'd5367, -32'd337},
{32'd6046, 32'd8773, 32'd573, -32'd11763},
{32'd3442, -32'd5582, -32'd14764, 32'd11912},
{-32'd1184, 32'd10686, -32'd4742, 32'd3647},
{-32'd6765, -32'd2341, 32'd3627, -32'd14256},
{32'd6671, 32'd13760, 32'd1695, 32'd3896},
{32'd468, -32'd1411, -32'd10781, -32'd4378},
{-32'd439, -32'd5456, 32'd4335, -32'd8601},
{32'd178, -32'd11978, -32'd13615, 32'd6177},
{32'd2917, -32'd8205, -32'd8575, 32'd7415},
{32'd5027, -32'd2203, -32'd348, 32'd425},
{32'd847, 32'd1068, 32'd3361, 32'd12445},
{-32'd2790, -32'd4217, -32'd12322, -32'd1998},
{32'd1044, -32'd4947, 32'd381, -32'd1889},
{32'd6414, 32'd5883, 32'd14080, 32'd5521},
{32'd8285, 32'd27441, 32'd2802, 32'd9369},
{-32'd5757, -32'd17536, 32'd1848, -32'd4862},
{-32'd6652, 32'd3594, 32'd758, -32'd4315},
{32'd14752, 32'd3861, 32'd4320, -32'd2321},
{-32'd5696, -32'd5541, -32'd4356, 32'd3504},
{32'd47, 32'd7581, 32'd944, -32'd9364},
{-32'd3390, 32'd253, -32'd6705, 32'd14975},
{-32'd10309, -32'd11324, 32'd8119, -32'd2076},
{-32'd17153, 32'd4365, -32'd33, 32'd1551},
{-32'd1134, -32'd5241, -32'd2291, 32'd12313},
{32'd4129, 32'd10061, -32'd5024, 32'd4069},
{-32'd5819, -32'd3069, 32'd903, -32'd9428},
{-32'd464, -32'd18200, -32'd662, 32'd5790},
{-32'd2838, -32'd6491, -32'd3784, 32'd3260},
{32'd1706, -32'd8034, -32'd711, -32'd5049},
{-32'd2022, 32'd1130, -32'd71, 32'd5066},
{32'd159, 32'd3644, -32'd958, 32'd841},
{32'd1142, 32'd13655, -32'd771, -32'd11476},
{-32'd11270, 32'd9827, -32'd4978, -32'd6996},
{32'd4353, 32'd1710, -32'd2400, 32'd2400},
{-32'd14966, 32'd9323, -32'd1145, 32'd2996},
{-32'd6547, 32'd4834, 32'd7845, 32'd8457},
{32'd8939, 32'd2820, 32'd2332, 32'd747},
{-32'd4192, -32'd2770, 32'd4281, -32'd2629},
{32'd15264, 32'd16172, 32'd10992, 32'd4267},
{-32'd1820, -32'd7280, -32'd1660, -32'd5486},
{-32'd6548, -32'd2597, -32'd6531, 32'd7928},
{-32'd5912, -32'd801, -32'd5106, 32'd5684},
{-32'd4304, 32'd17, 32'd5160, -32'd2568},
{32'd8879, 32'd18688, 32'd4339, -32'd6634},
{32'd1336, 32'd6820, 32'd3170, -32'd1784},
{-32'd4198, 32'd13422, -32'd897, -32'd8556},
{-32'd9261, -32'd813, -32'd2263, 32'd9242},
{32'd3471, 32'd1637, 32'd3913, -32'd861},
{-32'd1208, -32'd16331, -32'd4700, -32'd10296},
{-32'd9145, 32'd2619, -32'd2504, -32'd5225},
{-32'd8473, -32'd4047, 32'd460, 32'd5860},
{-32'd6369, 32'd8712, -32'd628, -32'd38},
{32'd12956, 32'd4416, 32'd1022, 32'd12630},
{-32'd8871, -32'd17969, -32'd10807, 32'd104},
{-32'd2372, -32'd58, -32'd8988, 32'd2102},
{-32'd272, -32'd4905, 32'd5995, 32'd2682},
{32'd294, -32'd7511, 32'd12295, 32'd5584},
{32'd3041, 32'd5703, 32'd9760, -32'd1422},
{32'd94, 32'd23454, 32'd174, -32'd2256},
{32'd7194, 32'd3527, 32'd1112, 32'd14628},
{32'd15890, 32'd9637, 32'd5196, 32'd3900},
{32'd1430, -32'd6105, -32'd1780, -32'd211},
{32'd5364, -32'd461, 32'd2998, 32'd9720},
{-32'd7102, 32'd8382, 32'd3920, 32'd3588},
{32'd8150, 32'd14279, 32'd6313, 32'd929},
{32'd11212, 32'd3343, -32'd10735, -32'd11453},
{-32'd5720, 32'd3997, -32'd5085, 32'd874},
{32'd6004, 32'd3915, 32'd5291, 32'd1343},
{32'd3478, -32'd18166, -32'd638, 32'd8224},
{32'd289, 32'd6346, -32'd3256, 32'd8255},
{32'd5587, 32'd1850, -32'd7037, -32'd3802},
{32'd4289, -32'd2605, -32'd6009, -32'd11830},
{32'd1460, 32'd2644, -32'd2474, -32'd5083},
{32'd8862, -32'd10696, -32'd4607, 32'd8699},
{-32'd2944, -32'd1047, -32'd6830, 32'd1392},
{32'd11635, -32'd3880, 32'd9908, 32'd1799},
{-32'd3331, -32'd18644, 32'd9472, 32'd7309},
{-32'd3933, 32'd5585, -32'd1223, 32'd6097},
{-32'd7300, -32'd7634, -32'd9542, -32'd727},
{32'd2645, 32'd17210, -32'd2572, -32'd5859},
{32'd2249, 32'd1357, 32'd5741, -32'd2563},
{-32'd15607, 32'd76, 32'd9764, 32'd3313},
{32'd6014, -32'd580, 32'd9665, -32'd6892},
{-32'd5696, 32'd2954, -32'd366, -32'd6344},
{-32'd7640, 32'd12026, -32'd1320, -32'd6203},
{32'd3993, 32'd778, 32'd5234, -32'd3891},
{-32'd4450, 32'd10644, 32'd6773, 32'd17860},
{32'd8566, 32'd2185, -32'd1962, 32'd5151},
{32'd1761, -32'd4494, -32'd5478, 32'd12641},
{-32'd2866, 32'd4552, 32'd4928, 32'd944},
{-32'd1133, -32'd7409, 32'd10859, 32'd10559},
{32'd11669, -32'd2701, -32'd4353, 32'd2015},
{-32'd4316, -32'd3786, 32'd9572, 32'd2812},
{32'd2330, -32'd3159, 32'd4682, 32'd5825},
{32'd19326, 32'd3547, -32'd1486, 32'd2956},
{-32'd2113, -32'd8516, -32'd7931, -32'd1364},
{-32'd4669, -32'd3014, -32'd1694, 32'd774},
{-32'd1524, -32'd1105, -32'd1052, -32'd8420},
{-32'd236, 32'd1459, 32'd4504, 32'd4723},
{-32'd12179, -32'd10416, -32'd10843, 32'd310},
{32'd11081, 32'd6155, -32'd3678, 32'd1264},
{-32'd1565, -32'd5244, -32'd4267, -32'd2807},
{-32'd3819, 32'd1470, 32'd9651, 32'd5448},
{32'd5869, 32'd3034, -32'd102, -32'd9222},
{-32'd17752, -32'd12317, -32'd3666, -32'd6928},
{32'd3305, 32'd10257, 32'd8819, -32'd11116},
{32'd1351, -32'd3079, -32'd3707, 32'd14077},
{-32'd8089, 32'd4572, 32'd5729, 32'd4239},
{32'd11448, -32'd3778, -32'd14994, -32'd3005},
{-32'd13573, -32'd12975, -32'd4290, -32'd8930},
{32'd6187, -32'd6321, -32'd11966, -32'd13178},
{32'd5690, 32'd14621, 32'd7366, 32'd422},
{32'd5338, -32'd6222, -32'd2461, -32'd4591},
{32'd5473, 32'd10834, 32'd4098, 32'd1465},
{-32'd7339, 32'd11897, -32'd4772, 32'd587},
{32'd10950, 32'd2485, 32'd1956, -32'd304},
{-32'd6427, -32'd2735, 32'd4842, -32'd161},
{32'd2001, -32'd4341, -32'd678, 32'd12282},
{-32'd7777, 32'd157, -32'd4215, -32'd3700},
{32'd1601, 32'd102, -32'd786, -32'd7731},
{-32'd6660, -32'd3911, -32'd355, 32'd4046},
{-32'd3463, 32'd2917, 32'd5975, -32'd3135},
{32'd24001, 32'd6414, 32'd1760, -32'd302},
{-32'd1138, 32'd1520, -32'd7971, -32'd3252},
{32'd11590, 32'd7838, 32'd6778, -32'd5342},
{32'd7970, 32'd7334, -32'd553, 32'd7655},
{32'd8370, -32'd70, -32'd1929, 32'd2577},
{32'd10783, 32'd5152, -32'd1812, -32'd7948},
{-32'd4959, 32'd1105, -32'd1337, 32'd3449},
{-32'd4898, 32'd8540, -32'd3724, -32'd8309},
{32'd9764, 32'd728, -32'd7464, -32'd791},
{-32'd9691, 32'd4371, -32'd684, -32'd9828},
{-32'd8597, -32'd487, -32'd8308, -32'd187},
{32'd13953, 32'd5878, 32'd6586, -32'd5876},
{-32'd4807, -32'd3057, 32'd472, -32'd1006},
{32'd5821, -32'd16340, 32'd6596, -32'd6317},
{32'd2701, 32'd2802, 32'd10804, 32'd3801},
{32'd2333, -32'd18312, -32'd1383, -32'd8908},
{-32'd2049, -32'd2099, 32'd6163, 32'd630},
{-32'd9893, -32'd10463, -32'd4777, -32'd1072},
{32'd12305, 32'd10761, -32'd1123, -32'd4067},
{-32'd7876, 32'd5376, -32'd4883, 32'd2128},
{-32'd286, 32'd2366, -32'd1899, -32'd394},
{-32'd2725, -32'd10354, -32'd175, 32'd5064},
{-32'd5162, -32'd5569, -32'd9527, -32'd7365},
{32'd7246, 32'd77, 32'd7762, -32'd12170},
{-32'd5643, -32'd5652, -32'd293, 32'd7241},
{32'd15956, -32'd300, 32'd11293, 32'd6380},
{32'd7683, -32'd2296, 32'd11559, 32'd2097},
{-32'd1670, 32'd1406, -32'd2770, -32'd14585},
{-32'd5453, -32'd2743, 32'd1650, 32'd3481},
{-32'd2052, -32'd8350, -32'd8131, 32'd6094},
{32'd6987, -32'd18822, 32'd5461, -32'd5699},
{-32'd12056, 32'd3923, 32'd7154, -32'd806},
{-32'd8736, -32'd3326, -32'd12414, -32'd2717},
{32'd4217, -32'd10264, 32'd872, -32'd1557},
{32'd3534, 32'd3551, 32'd1734, 32'd2525},
{-32'd7502, -32'd142, 32'd10905, 32'd9893},
{32'd8318, 32'd5867, 32'd1043, 32'd12343},
{32'd1517, 32'd2643, 32'd11808, 32'd990},
{-32'd5608, 32'd8814, 32'd7134, -32'd6110},
{32'd19513, 32'd16298, 32'd5114, -32'd6395},
{-32'd7305, -32'd3775, -32'd5215, -32'd346},
{-32'd10459, -32'd7274, 32'd243, -32'd7285},
{-32'd2709, -32'd19442, -32'd14476, 32'd9565},
{-32'd3392, 32'd1355, 32'd3101, 32'd1808},
{32'd2781, -32'd14102, -32'd6268, -32'd7669},
{32'd5155, -32'd4975, -32'd12889, 32'd1491},
{-32'd5743, 32'd330, 32'd4599, 32'd7544},
{32'd5172, 32'd8075, -32'd7932, -32'd10353},
{32'd19052, 32'd3778, -32'd5533, -32'd5851},
{32'd7541, 32'd6927, -32'd2389, -32'd2843},
{32'd5306, 32'd12077, -32'd966, -32'd1617},
{-32'd688, 32'd5681, 32'd1183, 32'd6713},
{-32'd3589, -32'd3937, -32'd1352, 32'd8174},
{32'd10934, -32'd8241, -32'd4257, 32'd4768},
{32'd9358, -32'd6048, 32'd1619, -32'd14632},
{32'd5437, -32'd799, 32'd5992, 32'd7115},
{32'd11342, 32'd4944, -32'd7758, 32'd2222},
{-32'd939, 32'd7089, -32'd4965, -32'd335},
{-32'd3652, -32'd4226, 32'd7633, 32'd6722},
{32'd794, -32'd615, -32'd3054, -32'd49},
{-32'd10125, -32'd9105, -32'd952, -32'd3690},
{32'd5731, 32'd15643, 32'd9639, -32'd9748},
{32'd3205, 32'd7540, 32'd10102, 32'd4819},
{32'd4360, -32'd8683, -32'd3831, 32'd3319},
{-32'd8176, -32'd248, 32'd5295, -32'd3530},
{-32'd7866, 32'd10577, -32'd3071, -32'd5493},
{-32'd8414, 32'd9224, 32'd5433, 32'd9909},
{32'd343, 32'd7174, 32'd811, -32'd3012},
{32'd407, 32'd8535, -32'd712, -32'd7242},
{32'd18546, 32'd6234, 32'd6929, 32'd3539},
{-32'd36, -32'd4585, -32'd161, 32'd1215},
{-32'd7165, 32'd550, -32'd5708, 32'd4231},
{-32'd13246, 32'd10404, -32'd2749, -32'd5975},
{-32'd6635, 32'd422, 32'd2890, -32'd1940},
{32'd526, -32'd536, 32'd4755, -32'd6742},
{32'd5392, -32'd8169, -32'd3216, 32'd4922},
{-32'd7254, -32'd1176, 32'd17936, 32'd7306},
{32'd530, -32'd5252, -32'd4418, -32'd6016},
{32'd1311, 32'd3356, -32'd9210, 32'd16452},
{-32'd2072, -32'd8486, -32'd4507, -32'd6244},
{32'd1575, -32'd7789, -32'd13462, -32'd4206},
{32'd16488, 32'd3772, 32'd327, -32'd9317},
{-32'd10106, 32'd3121, 32'd6188, 32'd4682},
{32'd486, -32'd6292, 32'd4991, 32'd2914},
{32'd1351, 32'd908, 32'd201, 32'd1486},
{-32'd2669, 32'd3704, -32'd5587, 32'd1962},
{-32'd10559, -32'd3259, -32'd8274, -32'd4808},
{32'd10398, -32'd5630, 32'd3126, 32'd2258},
{32'd3291, 32'd5343, 32'd4411, -32'd7692},
{-32'd4323, 32'd4412, 32'd13319, 32'd1591},
{32'd13742, -32'd7353, -32'd5450, -32'd4909},
{-32'd1505, -32'd1464, 32'd5614, 32'd11464},
{-32'd7158, 32'd3119, -32'd11168, -32'd4197},
{32'd6345, 32'd6985, 32'd8904, -32'd1545},
{32'd10643, 32'd3069, 32'd965, 32'd3770},
{-32'd1594, -32'd14057, -32'd689, 32'd4532},
{32'd9801, -32'd4237, -32'd2308, 32'd2720},
{32'd7938, 32'd13990, 32'd10361, -32'd1576},
{32'd11219, -32'd31, -32'd6344, -32'd4521},
{32'd3327, 32'd9038, 32'd10799, -32'd8130},
{-32'd6438, 32'd2417, -32'd7277, -32'd14841},
{-32'd3347, 32'd303, 32'd597, -32'd8000},
{-32'd12741, -32'd5130, -32'd12340, -32'd3216},
{-32'd1305, 32'd5865, -32'd468, -32'd511},
{-32'd246, -32'd7223, -32'd4983, -32'd7268},
{-32'd6911, 32'd16, 32'd3451, 32'd767},
{32'd1161, 32'd14079, -32'd16969, 32'd5769},
{32'd8394, 32'd2294, -32'd323, 32'd8162},
{32'd2104, 32'd5738, -32'd3446, -32'd1367},
{-32'd4478, -32'd8880, -32'd7857, -32'd4824},
{-32'd1521, -32'd503, 32'd1689, 32'd13798},
{32'd8315, -32'd2269, -32'd4860, -32'd2659},
{32'd4953, 32'd3298, 32'd1330, -32'd6124},
{-32'd17658, -32'd8109, -32'd7571, -32'd2033},
{-32'd11298, -32'd6714, -32'd1210, 32'd7727},
{-32'd1531, -32'd11064, 32'd7652, -32'd11230},
{-32'd317, 32'd16474, 32'd5999, -32'd2558}
},
{{32'd7054, -32'd1913, 32'd1886, 32'd6658},
{-32'd3585, 32'd2295, -32'd7767, 32'd248},
{32'd6593, -32'd3611, 32'd7072, -32'd1660},
{-32'd1145, 32'd3741, -32'd2918, 32'd7908},
{32'd9598, 32'd7151, -32'd6396, 32'd7101},
{-32'd2764, -32'd925, -32'd2980, 32'd1293},
{32'd4359, -32'd5042, -32'd677, 32'd1953},
{-32'd436, -32'd11694, -32'd5566, 32'd3736},
{32'd3055, -32'd6876, 32'd5752, -32'd1092},
{32'd3691, 32'd3955, 32'd2839, -32'd3201},
{-32'd15138, -32'd1432, 32'd361, 32'd12166},
{32'd5841, 32'd7860, -32'd1421, -32'd1630},
{32'd386, -32'd6628, -32'd3044, -32'd8871},
{32'd1636, 32'd366, 32'd3553, -32'd4386},
{32'd11305, 32'd118, 32'd3269, 32'd9891},
{-32'd11540, 32'd8881, -32'd738, 32'd533},
{32'd11881, 32'd1503, -32'd4133, -32'd3966},
{32'd4689, -32'd189, 32'd7477, -32'd9006},
{-32'd6603, 32'd4192, 32'd2860, 32'd9579},
{32'd491, 32'd10900, -32'd7025, 32'd4468},
{-32'd2337, 32'd1084, -32'd5381, 32'd5280},
{-32'd9234, 32'd305, -32'd1822, 32'd8254},
{-32'd2669, 32'd1170, -32'd4375, -32'd14546},
{-32'd10650, -32'd7759, 32'd4038, 32'd3053},
{32'd8421, 32'd4077, 32'd8553, -32'd1691},
{32'd4926, 32'd911, -32'd5773, -32'd3914},
{-32'd1771, -32'd6193, -32'd3089, -32'd7807},
{-32'd3706, -32'd3564, -32'd7270, -32'd9524},
{-32'd5518, 32'd15458, -32'd4466, 32'd13033},
{32'd9050, -32'd3500, 32'd6164, 32'd6664},
{-32'd879, -32'd1322, -32'd1801, -32'd2482},
{32'd478, 32'd389, -32'd2227, 32'd9060},
{32'd3348, -32'd1756, 32'd1516, 32'd1858},
{-32'd4988, 32'd8981, -32'd768, 32'd2231},
{32'd7669, 32'd3241, 32'd8768, 32'd2669},
{-32'd9327, 32'd3876, 32'd21807, 32'd5319},
{32'd5200, -32'd5368, 32'd187, -32'd136},
{32'd3266, 32'd11961, -32'd6175, 32'd3691},
{32'd917, 32'd1477, -32'd13173, -32'd6704},
{32'd4111, -32'd6508, 32'd3561, 32'd9330},
{-32'd15688, 32'd6271, 32'd755, 32'd207},
{-32'd6937, -32'd1559, 32'd11007, 32'd10398},
{32'd14102, 32'd12042, -32'd161, 32'd6071},
{32'd8677, 32'd1241, -32'd5435, -32'd4995},
{32'd2839, 32'd5621, 32'd3553, -32'd2038},
{-32'd5210, -32'd1658, -32'd8046, 32'd6742},
{-32'd6323, 32'd1075, 32'd5311, -32'd927},
{32'd109, 32'd5062, 32'd9663, 32'd1313},
{32'd2408, -32'd2589, 32'd1749, 32'd22},
{32'd6263, 32'd934, -32'd11417, -32'd4187},
{32'd6474, 32'd3430, 32'd262, -32'd9153},
{32'd851, 32'd5073, 32'd5526, 32'd2113},
{-32'd5003, 32'd1053, -32'd3115, 32'd12843},
{-32'd2322, 32'd5170, 32'd10317, 32'd424},
{32'd9585, -32'd3097, 32'd680, 32'd413},
{-32'd1528, 32'd3118, -32'd3997, -32'd4073},
{32'd6577, -32'd5872, -32'd13919, 32'd1752},
{-32'd971, -32'd1252, -32'd6706, 32'd8607},
{-32'd8676, 32'd3217, 32'd1922, 32'd4773},
{32'd6700, 32'd3583, -32'd2783, -32'd2494},
{-32'd1121, -32'd300, -32'd3522, 32'd8111},
{-32'd8610, -32'd12908, -32'd1371, 32'd1810},
{-32'd12157, -32'd1324, 32'd1472, 32'd1194},
{-32'd4066, 32'd1176, 32'd1703, 32'd1882},
{32'd7794, 32'd6742, -32'd11529, -32'd3753},
{32'd10884, -32'd2776, 32'd2127, 32'd3386},
{-32'd3113, -32'd387, -32'd10088, -32'd6804},
{32'd4329, -32'd6915, -32'd10844, -32'd5407},
{-32'd760, -32'd2683, -32'd4406, 32'd1029},
{-32'd2849, -32'd8644, 32'd15707, 32'd10259},
{32'd4132, -32'd232, -32'd7747, -32'd5715},
{32'd554, -32'd12717, -32'd1749, 32'd3928},
{-32'd1861, -32'd8502, 32'd5067, -32'd9623},
{-32'd6808, 32'd829, -32'd16746, 32'd9333},
{32'd9625, -32'd6629, -32'd7874, 32'd7124},
{32'd3432, -32'd8422, -32'd786, -32'd4642},
{-32'd1388, -32'd4301, 32'd2840, -32'd582},
{-32'd5810, -32'd1836, 32'd2420, 32'd2433},
{32'd3348, -32'd526, 32'd9837, -32'd10853},
{-32'd287, -32'd7508, -32'd1279, 32'd14146},
{32'd5530, 32'd3285, -32'd1468, -32'd13017},
{-32'd657, -32'd2029, 32'd1130, 32'd1513},
{-32'd8954, 32'd2677, -32'd2683, 32'd7556},
{-32'd12, 32'd15105, -32'd9972, -32'd7423},
{32'd12013, 32'd5537, 32'd4497, -32'd3109},
{-32'd7299, -32'd192, -32'd2520, 32'd4522},
{-32'd1485, 32'd8600, -32'd4893, 32'd4850},
{-32'd12659, -32'd298, 32'd4014, 32'd3724},
{-32'd4896, 32'd9556, -32'd5605, 32'd9321},
{32'd5289, 32'd7665, -32'd3918, -32'd1379},
{32'd107, 32'd1567, -32'd654, -32'd2826},
{32'd3081, -32'd3205, -32'd2805, 32'd4333},
{-32'd1791, -32'd1771, 32'd15371, -32'd1752},
{32'd8674, 32'd126, -32'd7553, -32'd5682},
{-32'd1854, -32'd2086, 32'd1026, -32'd6329},
{32'd7058, -32'd774, -32'd1305, -32'd6571},
{32'd3132, -32'd2463, -32'd1421, 32'd3027},
{32'd5496, -32'd97, 32'd13574, 32'd414},
{-32'd7266, -32'd2479, 32'd5174, 32'd123},
{32'd11680, 32'd429, 32'd1902, -32'd2062},
{32'd4125, -32'd2046, -32'd4315, -32'd2308},
{32'd4576, 32'd1056, 32'd8882, 32'd7006},
{-32'd5640, -32'd11742, -32'd2002, 32'd10416},
{-32'd11620, 32'd9346, -32'd5630, 32'd6453},
{32'd5112, 32'd2122, 32'd4470, 32'd3658},
{32'd4097, -32'd3942, -32'd1062, 32'd13523},
{-32'd7388, 32'd254, 32'd11840, -32'd7502},
{32'd4573, -32'd2564, 32'd458, -32'd2978},
{32'd11136, -32'd1435, 32'd7174, -32'd14791},
{32'd422, 32'd2014, -32'd2250, 32'd10671},
{-32'd5894, 32'd6583, -32'd50, -32'd2888},
{-32'd5700, -32'd1330, -32'd174, 32'd8042},
{-32'd3686, 32'd5586, -32'd8481, -32'd2117},
{32'd5196, -32'd1943, -32'd6623, -32'd9325},
{-32'd137, 32'd5492, 32'd1133, 32'd2598},
{32'd1098, 32'd1941, -32'd5253, -32'd3284},
{32'd2364, 32'd14915, 32'd3561, -32'd5741},
{32'd1402, -32'd2521, -32'd3057, -32'd8555},
{-32'd6753, 32'd334, -32'd2549, 32'd1911},
{32'd4102, 32'd447, -32'd103, 32'd1549},
{32'd7906, 32'd1499, -32'd3237, -32'd1439},
{32'd2471, -32'd5604, 32'd5463, 32'd9041},
{32'd4270, -32'd3180, -32'd10100, 32'd7459},
{-32'd2315, 32'd5683, -32'd2037, 32'd4862},
{32'd3420, -32'd2316, 32'd2006, 32'd12192},
{32'd10405, -32'd5666, -32'd14368, -32'd6634},
{32'd1203, 32'd1257, 32'd7982, -32'd5438},
{32'd2305, 32'd2454, -32'd2232, 32'd6717},
{-32'd7864, 32'd2425, -32'd3652, -32'd8140},
{-32'd10324, 32'd16955, 32'd7211, -32'd1725},
{-32'd483, 32'd8510, 32'd1407, 32'd5334},
{32'd474, -32'd3682, -32'd6358, 32'd599},
{-32'd6203, -32'd3610, -32'd1492, -32'd454},
{-32'd9724, -32'd10284, -32'd12563, -32'd761},
{32'd324, -32'd8370, -32'd1355, -32'd264},
{32'd1339, 32'd801, -32'd3342, -32'd8063},
{32'd1263, -32'd10909, -32'd253, 32'd11315},
{-32'd4028, 32'd10918, 32'd1027, -32'd3628},
{-32'd7162, 32'd4012, -32'd3220, -32'd8293},
{-32'd7139, -32'd2629, 32'd4612, -32'd8098},
{-32'd7907, -32'd2094, -32'd5637, -32'd6453},
{-32'd2798, -32'd3625, 32'd8320, -32'd379},
{32'd1605, 32'd4483, 32'd83, 32'd6019},
{32'd8799, 32'd3147, -32'd7223, 32'd6249},
{32'd7475, 32'd3161, 32'd2531, -32'd5588},
{32'd3044, -32'd8498, -32'd7864, -32'd5333},
{32'd5975, 32'd2094, -32'd3023, -32'd3742},
{-32'd1250, 32'd2841, 32'd6583, 32'd2687},
{32'd12924, -32'd5837, 32'd3401, 32'd6955},
{32'd719, 32'd405, 32'd3388, 32'd452},
{-32'd950, -32'd6716, 32'd3582, -32'd6767},
{-32'd5892, -32'd1404, 32'd94, 32'd3300},
{-32'd3558, -32'd1412, -32'd4452, -32'd30},
{-32'd369, -32'd8320, -32'd631, 32'd2246},
{-32'd1415, -32'd4041, 32'd4596, -32'd6270},
{32'd13081, -32'd2627, -32'd2055, 32'd3614},
{32'd4754, 32'd8001, 32'd18947, -32'd4581},
{32'd3291, 32'd11380, -32'd5274, 32'd2446},
{-32'd10456, 32'd1137, -32'd9330, 32'd12096},
{32'd2631, 32'd9785, 32'd13428, 32'd3699},
{-32'd13172, 32'd2322, 32'd1870, -32'd7145},
{32'd17071, -32'd2997, -32'd1944, -32'd1924},
{-32'd5310, 32'd3686, 32'd6621, 32'd16405},
{32'd9135, -32'd5662, -32'd1852, 32'd6596},
{32'd3051, 32'd2596, -32'd6405, 32'd7744},
{-32'd6193, 32'd4173, -32'd7339, 32'd3134},
{32'd4627, 32'd480, -32'd4543, -32'd8233},
{-32'd7106, 32'd135, -32'd8475, -32'd5198},
{-32'd3141, -32'd4485, -32'd151, 32'd2288},
{32'd10809, 32'd4666, 32'd5933, -32'd3278},
{-32'd10486, 32'd8146, 32'd8400, 32'd1015},
{32'd2165, -32'd1809, 32'd6249, 32'd8904},
{32'd1293, 32'd4174, 32'd3470, 32'd5131},
{-32'd9619, -32'd10678, -32'd31, 32'd2000},
{32'd8748, 32'd4362, 32'd7527, -32'd7096},
{-32'd2772, -32'd2048, 32'd5999, -32'd4775},
{32'd8960, 32'd1291, -32'd2724, -32'd2109},
{-32'd1835, 32'd11405, -32'd5615, -32'd2239},
{32'd1026, 32'd168, -32'd8900, 32'd5126},
{32'd5136, -32'd2862, -32'd7127, -32'd6946},
{32'd2280, 32'd3778, 32'd1792, -32'd2304},
{-32'd2603, 32'd4658, -32'd4914, 32'd8046},
{32'd152, -32'd1231, -32'd12232, 32'd634},
{-32'd1474, -32'd12012, 32'd62, 32'd11139},
{32'd8262, -32'd718, -32'd5529, -32'd11712},
{-32'd1243, 32'd8387, -32'd1335, -32'd4310},
{-32'd1940, -32'd6311, -32'd1130, 32'd1720},
{-32'd10810, -32'd13326, 32'd3212, 32'd3860},
{-32'd11114, 32'd27, -32'd5643, -32'd1262},
{-32'd2472, 32'd58, 32'd4353, 32'd1030},
{32'd10821, -32'd2217, 32'd7138, 32'd12118},
{32'd6262, -32'd638, 32'd6868, 32'd5640},
{-32'd804, 32'd5196, -32'd6137, -32'd4780},
{-32'd11334, -32'd3883, 32'd6899, 32'd24},
{-32'd5407, 32'd6759, -32'd10054, -32'd14663},
{32'd8343, 32'd10249, 32'd4289, -32'd3145},
{32'd3510, 32'd7030, 32'd5180, -32'd6542},
{-32'd695, -32'd273, -32'd1328, -32'd701},
{-32'd1723, -32'd6423, 32'd3569, -32'd8974},
{32'd4968, -32'd83, 32'd1651, -32'd3541},
{-32'd1956, -32'd2531, -32'd564, -32'd1551},
{32'd448, -32'd10481, -32'd441, -32'd8049},
{-32'd8373, -32'd11134, -32'd10263, 32'd3972},
{-32'd8629, -32'd9264, -32'd8864, 32'd9043},
{-32'd2969, 32'd4836, -32'd1787, 32'd5930},
{-32'd4180, 32'd4044, -32'd2628, 32'd7801},
{32'd787, 32'd2733, -32'd4043, -32'd2747},
{-32'd2284, 32'd3378, -32'd1336, 32'd1234},
{32'd9901, -32'd7705, -32'd1287, -32'd2646},
{32'd282, 32'd776, -32'd576, 32'd3390},
{-32'd10544, -32'd7180, -32'd685, -32'd12002},
{32'd1102, 32'd10290, -32'd4833, -32'd6301},
{-32'd13041, 32'd185, -32'd8557, 32'd4516},
{32'd1551, 32'd10426, 32'd8436, 32'd511},
{32'd11457, -32'd8814, -32'd1675, -32'd823},
{32'd3295, 32'd1330, 32'd7352, 32'd8991},
{-32'd8994, 32'd4443, -32'd3708, -32'd1751},
{-32'd3287, -32'd2231, -32'd4235, -32'd13777},
{32'd8200, -32'd2951, -32'd4067, 32'd1820},
{32'd4673, -32'd13040, 32'd1901, 32'd1201},
{32'd4145, -32'd5841, -32'd11483, -32'd649},
{-32'd1609, 32'd1261, 32'd72, 32'd3217},
{32'd13904, -32'd1976, 32'd417, 32'd3641},
{-32'd2963, 32'd1589, 32'd3486, -32'd4801},
{32'd2450, 32'd1813, 32'd4167, -32'd2107},
{-32'd8341, 32'd7854, -32'd5863, 32'd10306},
{-32'd1846, 32'd5936, -32'd3946, 32'd3901},
{-32'd6072, 32'd861, -32'd475, -32'd8011},
{-32'd2503, 32'd12162, 32'd5012, 32'd10421},
{32'd1077, -32'd3037, 32'd645, 32'd7964},
{32'd736, -32'd9815, 32'd4292, -32'd3002},
{-32'd7521, 32'd5479, -32'd3924, 32'd11569},
{-32'd4035, 32'd1783, 32'd12136, -32'd2504},
{32'd4011, -32'd11290, -32'd70, -32'd11095},
{32'd645, -32'd2098, -32'd1037, -32'd8617},
{-32'd10328, -32'd7534, -32'd4676, -32'd4741},
{32'd4307, 32'd1966, -32'd8568, 32'd505},
{-32'd5599, -32'd9037, -32'd8128, -32'd3492},
{32'd10563, -32'd2337, 32'd1623, 32'd1612},
{-32'd6113, -32'd10952, 32'd1901, 32'd5979},
{-32'd3640, -32'd3052, 32'd171, 32'd5377},
{-32'd5347, -32'd8890, -32'd6865, 32'd3459},
{-32'd107, 32'd53, -32'd8692, 32'd2016},
{-32'd3080, 32'd6010, -32'd16107, -32'd5574},
{32'd3883, 32'd5077, 32'd3693, 32'd3648},
{32'd4415, -32'd4650, 32'd9851, -32'd4131},
{32'd2582, -32'd6100, 32'd10961, -32'd3163},
{32'd2238, 32'd3045, 32'd8626, -32'd5278},
{32'd9156, -32'd1770, 32'd10214, 32'd4625},
{32'd1373, -32'd632, -32'd6563, -32'd5475},
{-32'd2680, 32'd393, -32'd1816, -32'd6628},
{32'd10089, -32'd1322, 32'd6649, 32'd3177},
{32'd12895, 32'd5144, -32'd6550, -32'd4953},
{-32'd232, 32'd1944, -32'd87, 32'd455},
{-32'd5884, -32'd1247, -32'd1238, 32'd5359},
{-32'd1566, 32'd6967, 32'd2230, 32'd5270},
{-32'd7115, 32'd5766, -32'd5794, -32'd4713},
{32'd2307, -32'd3647, -32'd5122, -32'd3001},
{-32'd12070, -32'd1219, -32'd39, 32'd7124},
{32'd4510, -32'd5274, -32'd5957, 32'd7430},
{-32'd623, 32'd10578, -32'd2376, -32'd2731},
{32'd9644, 32'd2776, 32'd12445, 32'd848},
{32'd12734, 32'd7862, 32'd4792, -32'd13706},
{-32'd1414, -32'd6714, -32'd4456, 32'd6640},
{32'd3962, -32'd1566, -32'd4615, -32'd5109},
{-32'd1211, 32'd2412, 32'd5226, 32'd5590},
{32'd9798, -32'd664, 32'd2325, -32'd1198},
{-32'd3370, 32'd10149, 32'd7226, -32'd237},
{32'd3923, 32'd1637, 32'd375, 32'd11443},
{32'd3171, -32'd146, 32'd1219, -32'd11161},
{-32'd2558, 32'd6178, -32'd1531, 32'd9827},
{32'd2414, 32'd2322, -32'd7643, -32'd10174},
{-32'd1148, 32'd5823, 32'd1237, 32'd732},
{-32'd3906, 32'd1881, 32'd4306, -32'd4431},
{32'd5031, 32'd1797, -32'd5438, -32'd7396},
{-32'd11651, -32'd503, 32'd8645, 32'd6941},
{32'd5076, 32'd3396, 32'd4686, 32'd3131},
{32'd4397, -32'd53, -32'd2107, -32'd2735},
{-32'd2270, 32'd690, -32'd1700, -32'd309},
{32'd1632, -32'd7833, -32'd1915, 32'd3776},
{-32'd796, 32'd95, 32'd8168, 32'd2474},
{-32'd2320, -32'd2381, -32'd13522, 32'd5976},
{32'd11876, -32'd3450, -32'd7102, -32'd2564},
{-32'd7644, -32'd3211, 32'd5072, 32'd1763},
{32'd33, 32'd11822, -32'd1318, -32'd2620},
{-32'd11941, -32'd2854, -32'd2821, -32'd4030},
{32'd1491, -32'd848, -32'd11692, -32'd2535},
{-32'd5124, -32'd10203, 32'd2508, -32'd7645},
{-32'd6070, -32'd2978, 32'd8684, -32'd6485},
{32'd5658, 32'd4065, 32'd3592, 32'd12352},
{-32'd6064, -32'd2988, 32'd1011, 32'd18},
{32'd4697, 32'd370, 32'd1081, 32'd5343},
{-32'd848, 32'd5586, -32'd2014, 32'd8517},
{-32'd848, 32'd686, 32'd2298, 32'd918},
{-32'd4780, -32'd174, 32'd7016, -32'd3134},
{32'd6575, -32'd7407, 32'd7291, 32'd248},
{-32'd595, -32'd4812, 32'd5770, 32'd316},
{-32'd2437, 32'd9517, 32'd8787, 32'd11370},
{32'd10731, 32'd864, 32'd1101, 32'd3293},
{-32'd9095, 32'd968, 32'd3254, 32'd1790}
},
{{-32'd222, 32'd2196, -32'd4194, -32'd4},
{-32'd1274, -32'd11517, -32'd4344, 32'd1118},
{32'd1297, 32'd12849, -32'd1250, 32'd5432},
{-32'd2112, 32'd7009, 32'd10789, -32'd6169},
{32'd8563, 32'd11219, 32'd3777, -32'd1725},
{-32'd4137, -32'd992, 32'd16185, -32'd7746},
{32'd3071, -32'd4854, 32'd8653, -32'd6222},
{-32'd9083, -32'd21221, 32'd8711, -32'd388},
{-32'd2113, -32'd1691, 32'd7585, -32'd2024},
{-32'd3330, -32'd2144, -32'd845, 32'd732},
{32'd8073, 32'd9009, 32'd6403, 32'd1190},
{-32'd8836, -32'd13839, 32'd1732, -32'd2422},
{32'd3974, 32'd4670, 32'd2708, -32'd11012},
{32'd5746, 32'd1084, -32'd2562, -32'd2944},
{32'd2974, 32'd7752, -32'd5786, -32'd4644},
{-32'd5449, 32'd977, -32'd7571, 32'd3194},
{-32'd7227, 32'd7385, -32'd5915, -32'd5802},
{32'd13639, 32'd12253, -32'd5083, 32'd5066},
{32'd2310, -32'd13272, -32'd10786, -32'd11839},
{-32'd9566, -32'd13842, 32'd3216, 32'd229},
{32'd7150, 32'd6138, 32'd7306, -32'd15239},
{32'd8175, 32'd14589, -32'd2383, -32'd1905},
{-32'd2011, 32'd6744, -32'd10889, -32'd9245},
{32'd54, 32'd3544, -32'd7605, 32'd5527},
{32'd4983, -32'd13314, 32'd5923, 32'd530},
{32'd155, 32'd2990, -32'd938, -32'd2771},
{-32'd4362, -32'd8057, -32'd7215, -32'd4392},
{-32'd5842, 32'd12787, -32'd1922, -32'd5999},
{-32'd4048, 32'd8573, -32'd639, -32'd15352},
{32'd9119, 32'd7989, 32'd3564, 32'd13046},
{32'd3248, 32'd10168, 32'd2359, -32'd2344},
{32'd3988, 32'd5124, -32'd2260, -32'd1824},
{32'd1057, -32'd8399, -32'd2291, 32'd6694},
{-32'd3295, 32'd2526, -32'd6645, 32'd2209},
{32'd431, -32'd4389, 32'd4566, 32'd3646},
{32'd5220, -32'd9428, 32'd5324, 32'd12490},
{-32'd4351, 32'd7956, -32'd14971, 32'd7285},
{32'd5969, -32'd3256, -32'd4592, -32'd1128},
{-32'd7160, 32'd3523, -32'd10212, 32'd1450},
{-32'd876, -32'd17443, -32'd8773, 32'd11901},
{32'd6786, -32'd10555, -32'd3749, -32'd3435},
{32'd9067, -32'd7259, 32'd13808, -32'd2907},
{-32'd493, -32'd5628, 32'd5698, 32'd9996},
{-32'd2969, -32'd4788, -32'd12797, -32'd3561},
{-32'd10071, -32'd14862, -32'd7005, 32'd9415},
{-32'd5164, 32'd12536, -32'd6441, 32'd4693},
{-32'd589, -32'd14930, 32'd8457, 32'd1720},
{32'd3206, -32'd1513, -32'd8428, -32'd12106},
{-32'd5288, -32'd8267, 32'd7084, -32'd4918},
{-32'd1664, -32'd5863, 32'd1343, 32'd3495},
{-32'd3442, 32'd7614, 32'd6794, -32'd13590},
{32'd2457, -32'd13532, -32'd1193, 32'd8149},
{32'd776, -32'd237, -32'd8894, -32'd14060},
{32'd7222, -32'd4650, -32'd10075, -32'd4061},
{32'd6644, 32'd7030, -32'd10684, 32'd4895},
{-32'd2397, 32'd1300, 32'd12265, 32'd2284},
{-32'd2157, 32'd18892, -32'd1531, -32'd620},
{32'd3442, 32'd11420, -32'd5380, 32'd1891},
{-32'd1420, -32'd1754, -32'd8167, -32'd1050},
{-32'd16636, -32'd765, 32'd15368, 32'd1684},
{32'd3461, 32'd11233, 32'd4631, 32'd2213},
{32'd9435, -32'd10658, -32'd2953, -32'd10861},
{32'd1982, -32'd564, -32'd9105, -32'd1122},
{-32'd6748, 32'd6339, -32'd2928, -32'd4929},
{-32'd5360, -32'd680, -32'd4809, 32'd11442},
{32'd103, -32'd2612, 32'd11225, -32'd5518},
{32'd888, -32'd3131, -32'd2456, -32'd3948},
{-32'd5064, 32'd5953, -32'd505, -32'd3492},
{-32'd3046, -32'd16181, -32'd19472, -32'd5693},
{-32'd10841, -32'd5000, 32'd4128, 32'd2268},
{-32'd3981, 32'd5629, -32'd3730, 32'd11350},
{-32'd158, 32'd1181, 32'd12062, 32'd7544},
{32'd9981, -32'd811, -32'd6073, 32'd2686},
{-32'd7632, 32'd15308, 32'd1303, -32'd4870},
{-32'd2531, 32'd12004, 32'd8810, 32'd1419},
{32'd5829, -32'd4298, -32'd3516, 32'd18841},
{32'd335, -32'd7995, -32'd4676, -32'd3979},
{32'd4074, 32'd2826, 32'd4284, -32'd2441},
{-32'd5304, -32'd2140, 32'd13868, -32'd12174},
{32'd2836, 32'd2195, -32'd13401, 32'd13918},
{-32'd4941, -32'd15881, -32'd3281, -32'd19931},
{32'd2576, 32'd1451, -32'd4991, -32'd7622},
{-32'd5091, 32'd17487, 32'd2484, 32'd7609},
{32'd3823, -32'd1147, 32'd12559, 32'd5078},
{32'd11402, -32'd6614, 32'd12452, 32'd12678},
{32'd1306, 32'd20199, 32'd969, 32'd651},
{-32'd71, 32'd1462, -32'd11153, 32'd7958},
{32'd1201, 32'd5322, -32'd14102, 32'd435},
{-32'd14392, 32'd5201, 32'd6516, 32'd4868},
{-32'd9467, 32'd7973, 32'd5270, 32'd9531},
{-32'd6468, -32'd1714, -32'd7, 32'd937},
{32'd2568, 32'd2373, -32'd1709, 32'd609},
{32'd2117, -32'd14685, -32'd1055, -32'd11946},
{-32'd2216, 32'd12042, 32'd3411, -32'd3348},
{32'd2973, 32'd898, 32'd2335, 32'd15433},
{32'd3940, -32'd20722, -32'd5337, -32'd14480},
{-32'd1023, 32'd2093, -32'd2799, 32'd6204},
{32'd4422, -32'd102, 32'd284, 32'd14037},
{-32'd2524, 32'd15227, 32'd8295, -32'd205},
{32'd3344, 32'd5207, -32'd1246, 32'd158},
{32'd5013, 32'd316, -32'd16160, -32'd4408},
{-32'd1319, -32'd3784, 32'd4037, 32'd3350},
{-32'd4665, 32'd5350, -32'd6456, 32'd9057},
{-32'd191, 32'd3200, 32'd236, -32'd13936},
{-32'd745, 32'd2503, -32'd5587, -32'd2486},
{32'd15021, -32'd3708, -32'd1569, 32'd4228},
{32'd4160, 32'd10589, 32'd12478, -32'd4823},
{32'd1231, 32'd1515, -32'd6384, -32'd3398},
{32'd2505, 32'd4162, -32'd10028, -32'd16564},
{-32'd3501, 32'd6835, -32'd5785, 32'd2339},
{-32'd5316, 32'd9629, -32'd7247, -32'd6111},
{-32'd2305, -32'd7095, -32'd17525, 32'd3248},
{-32'd11944, 32'd3531, -32'd17767, 32'd4580},
{32'd8592, -32'd2982, 32'd5527, 32'd6854},
{32'd3177, -32'd12455, -32'd3369, -32'd1568},
{-32'd5279, -32'd1830, 32'd2618, -32'd5650},
{-32'd1288, -32'd979, 32'd10897, -32'd6007},
{-32'd2817, -32'd6233, 32'd12238, -32'd2927},
{-32'd7937, 32'd19856, 32'd10417, -32'd7847},
{-32'd5362, -32'd4006, 32'd4762, 32'd6657},
{-32'd6986, -32'd2712, -32'd9222, -32'd4782},
{32'd5833, -32'd3474, -32'd4525, 32'd9779},
{-32'd5800, -32'd4486, 32'd1628, -32'd6742},
{32'd6194, 32'd5038, 32'd14098, -32'd603},
{32'd4385, -32'd5463, 32'd1430, 32'd10814},
{-32'd9184, -32'd2532, 32'd38, 32'd7847},
{32'd9515, -32'd21459, 32'd9201, -32'd3751},
{-32'd1321, 32'd12545, -32'd1414, 32'd5320},
{32'd6518, -32'd9418, -32'd5104, -32'd6754},
{-32'd8040, -32'd16259, -32'd4711, 32'd6016},
{32'd9607, 32'd3105, 32'd790, 32'd4217},
{-32'd1686, -32'd27276, -32'd83, 32'd1655},
{32'd3081, -32'd15078, -32'd7915, -32'd17161},
{-32'd2979, -32'd1356, 32'd4818, -32'd13108},
{-32'd3582, -32'd4843, -32'd7495, 32'd1474},
{-32'd8380, -32'd8014, 32'd13268, 32'd4928},
{-32'd4329, 32'd2249, 32'd7939, 32'd11359},
{-32'd6577, -32'd11027, -32'd14168, 32'd7758},
{32'd7807, -32'd2243, 32'd6634, -32'd1480},
{-32'd8027, -32'd12354, -32'd11387, -32'd18882},
{-32'd3247, -32'd339, -32'd14135, -32'd2679},
{32'd3282, 32'd2563, 32'd2398, 32'd3876},
{32'd2341, 32'd7941, 32'd5656, 32'd2253},
{32'd1289, 32'd11109, 32'd5494, -32'd15276},
{32'd7663, 32'd169, -32'd4935, 32'd496},
{-32'd1040, 32'd16363, -32'd1595, 32'd3326},
{32'd2552, -32'd5777, -32'd13850, 32'd0},
{32'd926, -32'd1201, 32'd4017, -32'd1507},
{-32'd4610, -32'd7644, 32'd13575, -32'd9938},
{-32'd7068, -32'd11451, 32'd5776, -32'd2343},
{32'd4754, 32'd70, -32'd9146, 32'd9752},
{-32'd6898, -32'd8710, 32'd10054, -32'd6043},
{32'd107, 32'd6720, -32'd11819, -32'd1663},
{-32'd4729, 32'd8380, 32'd3702, 32'd2288},
{-32'd3133, -32'd4490, 32'd2852, 32'd3031},
{-32'd4436, 32'd2691, -32'd7112, 32'd6900},
{-32'd8444, -32'd6639, 32'd9638, 32'd8114},
{-32'd5016, 32'd2694, 32'd4267, 32'd1274},
{32'd3295, 32'd5350, -32'd16890, -32'd578},
{-32'd166, -32'd8966, 32'd11536, 32'd8861},
{-32'd4339, 32'd9018, -32'd462, -32'd7167},
{-32'd895, -32'd15630, 32'd7967, 32'd5903},
{-32'd5, 32'd3871, -32'd9795, -32'd15593},
{32'd1526, 32'd9491, -32'd223, -32'd4877},
{-32'd8950, -32'd3336, 32'd2174, 32'd7758},
{-32'd11839, 32'd9283, 32'd568, 32'd2863},
{32'd10713, -32'd1495, 32'd1355, -32'd4659},
{-32'd6653, -32'd8666, 32'd3447, 32'd14993},
{32'd10729, -32'd704, -32'd11654, 32'd8899},
{32'd13318, -32'd3711, -32'd4419, 32'd6270},
{32'd4157, -32'd1395, 32'd9983, -32'd9321},
{32'd2094, -32'd15055, 32'd14696, -32'd2519},
{-32'd5555, -32'd6258, 32'd4609, 32'd3350},
{32'd6253, -32'd5984, -32'd4215, -32'd11364},
{32'd726, 32'd5850, 32'd14832, -32'd6127},
{32'd5775, -32'd7610, -32'd11936, 32'd1075},
{-32'd2006, -32'd8641, -32'd6574, 32'd8421},
{-32'd11495, 32'd4749, 32'd1239, -32'd4780},
{32'd860, -32'd1929, -32'd11208, 32'd7333},
{-32'd534, 32'd14026, -32'd979, -32'd7438},
{-32'd1114, -32'd8619, -32'd8230, 32'd7917},
{-32'd1408, -32'd1366, -32'd21353, 32'd8665},
{32'd1029, -32'd9352, 32'd1175, -32'd1367},
{-32'd1245, -32'd11428, 32'd9459, 32'd9198},
{-32'd1964, 32'd6131, -32'd8244, 32'd3390},
{-32'd512, -32'd8578, 32'd17296, -32'd13831},
{-32'd7167, -32'd4162, 32'd16270, -32'd6037},
{-32'd2111, 32'd13350, -32'd7812, 32'd7987},
{-32'd10681, 32'd17047, 32'd9193, 32'd1328},
{32'd6197, 32'd13679, -32'd94, 32'd2546},
{32'd5050, -32'd15764, 32'd4611, 32'd57},
{-32'd1008, -32'd1490, -32'd15356, -32'd6030},
{32'd4275, 32'd14588, -32'd1859, 32'd1656},
{32'd1277, -32'd3547, -32'd968, -32'd9477},
{-32'd7145, 32'd885, 32'd4679, 32'd7891},
{-32'd614, -32'd23537, -32'd18038, 32'd3253},
{32'd13581, -32'd16692, -32'd8093, -32'd1361},
{32'd1366, 32'd5966, -32'd356, 32'd7706},
{-32'd7876, 32'd4975, 32'd14874, -32'd12752},
{32'd3169, -32'd25939, -32'd4460, 32'd1850},
{32'd172, -32'd2409, -32'd2067, -32'd1991},
{-32'd2624, -32'd11596, 32'd1722, -32'd2174},
{-32'd6868, 32'd2258, -32'd5407, -32'd5207},
{-32'd1331, 32'd7785, 32'd544, -32'd8548},
{-32'd7335, 32'd2579, 32'd2431, 32'd2927},
{32'd10582, 32'd3609, 32'd6360, 32'd306},
{32'd7087, 32'd9665, 32'd7321, 32'd1525},
{-32'd12009, 32'd497, 32'd6838, -32'd9485},
{-32'd314, 32'd5997, 32'd483, 32'd1090},
{32'd2168, -32'd10787, 32'd2761, 32'd15287},
{32'd1755, 32'd5203, 32'd3811, 32'd2114},
{-32'd8324, -32'd7768, -32'd499, 32'd2003},
{32'd4323, 32'd6963, 32'd4107, 32'd12270},
{-32'd234, -32'd9582, -32'd5034, -32'd1870},
{-32'd9668, -32'd5001, -32'd17249, -32'd5608},
{32'd10733, 32'd5814, -32'd4418, -32'd14957},
{-32'd11330, 32'd5634, 32'd26096, 32'd9511},
{-32'd4427, 32'd19686, 32'd4453, -32'd8407},
{-32'd453, 32'd9209, 32'd3681, 32'd11168},
{32'd6525, 32'd4425, 32'd10453, -32'd1588},
{-32'd4059, 32'd22603, 32'd4187, 32'd7025},
{32'd5646, 32'd6008, -32'd7372, -32'd6070},
{-32'd9001, 32'd13941, -32'd3507, -32'd1019},
{32'd11202, 32'd7261, -32'd2060, 32'd4319},
{32'd3497, 32'd14630, -32'd2420, -32'd9098},
{-32'd9402, 32'd10826, -32'd1877, 32'd17845},
{32'd5267, 32'd4999, 32'd12556, -32'd9182},
{32'd2919, -32'd12696, -32'd1215, -32'd205},
{32'd1201, -32'd12344, 32'd1439, -32'd9761},
{-32'd8322, 32'd4975, 32'd9178, 32'd7252},
{32'd6305, -32'd4680, -32'd3489, -32'd262},
{32'd1161, -32'd7021, -32'd7500, -32'd4204},
{32'd5481, 32'd7129, 32'd8567, 32'd3311},
{-32'd950, 32'd3845, -32'd2836, 32'd6225},
{32'd1402, -32'd8401, 32'd8768, 32'd11931},
{-32'd2090, 32'd5108, -32'd3530, 32'd15496},
{32'd9204, 32'd1905, -32'd299, -32'd8486},
{32'd7928, 32'd5599, -32'd7985, 32'd1273},
{32'd6358, 32'd3442, 32'd1616, -32'd204},
{32'd2677, -32'd5814, 32'd1154, 32'd8224},
{32'd2421, 32'd1030, -32'd6270, 32'd10093},
{-32'd240, 32'd5995, 32'd8671, 32'd1231},
{32'd1856, 32'd5795, 32'd2368, -32'd190},
{-32'd11183, 32'd12365, 32'd2443, 32'd4170},
{-32'd1861, 32'd4836, -32'd4386, 32'd2633},
{32'd15280, -32'd3340, -32'd5420, 32'd4078},
{32'd7528, -32'd6967, 32'd12184, -32'd4704},
{32'd6739, -32'd15462, 32'd13445, -32'd3144},
{32'd14713, 32'd11491, 32'd13377, -32'd1414},
{-32'd1022, 32'd16370, 32'd480, 32'd3536},
{-32'd1746, 32'd3511, 32'd10418, -32'd14242},
{32'd4448, -32'd12198, -32'd21238, -32'd14154},
{-32'd4739, 32'd7113, -32'd15146, 32'd4719},
{32'd10308, 32'd13828, -32'd2410, -32'd18567},
{32'd3404, 32'd12198, -32'd5852, -32'd1611},
{-32'd560, 32'd11907, -32'd4036, -32'd4568},
{-32'd3480, -32'd12516, 32'd1823, -32'd4715},
{-32'd11524, 32'd10796, -32'd4972, 32'd945},
{32'd3397, -32'd4429, -32'd13638, 32'd3740},
{32'd4511, 32'd1696, 32'd2675, 32'd12224},
{32'd1271, -32'd3000, 32'd13286, 32'd10058},
{32'd14162, 32'd7260, 32'd7066, 32'd8458},
{32'd6575, -32'd4779, 32'd1441, 32'd4641},
{32'd4796, -32'd8788, -32'd8424, -32'd9991},
{-32'd2348, -32'd6973, 32'd7563, -32'd5556},
{-32'd705, 32'd481, 32'd6401, -32'd3221},
{32'd2990, 32'd5426, -32'd1666, 32'd5545},
{32'd3077, -32'd2724, -32'd12259, 32'd4999},
{32'd4060, -32'd7974, 32'd3636, 32'd6544},
{-32'd2876, 32'd5088, 32'd2445, 32'd14559},
{32'd1283, 32'd10095, 32'd6149, -32'd4797},
{-32'd1985, 32'd11511, 32'd3379, -32'd1400},
{32'd6429, 32'd576, 32'd315, -32'd6357},
{32'd11866, -32'd3930, 32'd6503, 32'd3684},
{32'd24255, 32'd3312, 32'd556, -32'd7962},
{32'd12316, -32'd240, -32'd3623, 32'd5048},
{32'd2614, 32'd1583, -32'd1913, 32'd4579},
{-32'd2200, -32'd6869, 32'd2401, -32'd18815},
{32'd3909, 32'd3368, -32'd1203, 32'd1042},
{-32'd2385, -32'd7368, -32'd9046, 32'd6868},
{-32'd6603, 32'd158, 32'd2849, 32'd5401},
{-32'd17026, 32'd6791, 32'd3659, 32'd7515},
{-32'd5894, 32'd16802, 32'd3231, -32'd2562},
{-32'd609, 32'd3751, 32'd19586, -32'd6196},
{-32'd11264, -32'd2320, -32'd6858, 32'd4208},
{-32'd11935, -32'd15205, -32'd851, -32'd8382},
{-32'd12807, 32'd11327, 32'd5307, -32'd6666},
{32'd4764, -32'd1769, -32'd5506, 32'd9106},
{32'd9054, -32'd2748, 32'd2758, -32'd5963},
{32'd7686, -32'd10042, -32'd15554, 32'd4027},
{-32'd6311, 32'd12487, -32'd5480, -32'd2868},
{-32'd4830, -32'd9509, 32'd1860, 32'd6732},
{32'd1935, 32'd847, -32'd2925, -32'd6700},
{32'd2293, -32'd7569, 32'd2918, -32'd1654},
{-32'd2074, -32'd3810, 32'd2427, -32'd7163},
{32'd13290, -32'd5230, -32'd1876, 32'd5716},
{32'd2140, -32'd7847, -32'd11608, 32'd3175},
{32'd5363, -32'd3876, 32'd2453, 32'd403},
{-32'd10180, -32'd7248, 32'd7778, -32'd6110},
{-32'd7783, -32'd10046, -32'd16118, 32'd11065}
},
{{-32'd3084, 32'd14766, 32'd10686, 32'd1042},
{-32'd8029, -32'd8046, -32'd11608, -32'd12397},
{-32'd8925, 32'd2236, 32'd3199, 32'd12851},
{32'd350, 32'd5765, 32'd7064, -32'd1433},
{32'd9676, -32'd11017, -32'd1007, 32'd1698},
{-32'd8508, -32'd11439, -32'd10803, -32'd2850},
{32'd3302, -32'd11136, 32'd5733, 32'd8146},
{32'd12053, -32'd1569, -32'd5981, 32'd3344},
{-32'd29, -32'd11184, -32'd14361, -32'd2063},
{32'd584, 32'd7625, 32'd12049, 32'd3619},
{32'd1965, -32'd3770, -32'd1225, -32'd17117},
{-32'd19945, 32'd7632, -32'd1076, -32'd11725},
{32'd3029, -32'd7120, -32'd5228, -32'd3697},
{32'd2821, -32'd2929, 32'd8201, 32'd1816},
{32'd10532, -32'd12179, -32'd6132, -32'd1760},
{32'd6321, -32'd1825, -32'd3913, 32'd319},
{32'd6533, 32'd14028, 32'd5140, 32'd3128},
{32'd2912, 32'd2660, 32'd7108, 32'd3320},
{32'd15673, -32'd3060, -32'd3230, -32'd1646},
{32'd4703, 32'd6904, 32'd3186, 32'd3125},
{32'd3155, 32'd4735, 32'd13021, 32'd5887},
{-32'd1847, -32'd7432, -32'd3318, -32'd2757},
{32'd8867, -32'd6526, -32'd8463, 32'd3190},
{32'd189, -32'd2156, -32'd10655, 32'd12869},
{32'd13495, 32'd784, 32'd9476, 32'd7469},
{-32'd2882, 32'd3137, 32'd1482, 32'd12090},
{-32'd10905, -32'd21644, 32'd3004, -32'd7925},
{32'd7068, 32'd10568, -32'd2008, 32'd594},
{-32'd12613, 32'd5452, 32'd23916, -32'd7061},
{32'd1291, -32'd14125, -32'd3442, -32'd363},
{-32'd2696, -32'd16517, -32'd13877, 32'd13799},
{-32'd3844, -32'd12071, -32'd2710, 32'd3391},
{32'd1700, 32'd17263, -32'd5492, -32'd2093},
{32'd1223, 32'd3439, -32'd8519, 32'd3073},
{32'd4900, -32'd1445, 32'd2523, 32'd1138},
{32'd3490, 32'd5714, -32'd8742, -32'd7914},
{32'd4629, -32'd2194, 32'd6693, 32'd13537},
{-32'd120, 32'd41, 32'd6629, 32'd87},
{-32'd10192, 32'd372, 32'd2599, -32'd9325},
{-32'd12419, 32'd5166, -32'd11170, -32'd4291},
{32'd1038, 32'd1329, -32'd1143, 32'd3091},
{32'd493, 32'd2205, -32'd3969, -32'd4892},
{-32'd9040, 32'd8208, 32'd309, -32'd6636},
{32'd2045, 32'd8432, -32'd6742, -32'd149},
{32'd1047, 32'd13051, -32'd12151, 32'd11811},
{-32'd10136, 32'd5501, -32'd2503, -32'd10999},
{32'd10853, 32'd5646, -32'd7690, -32'd700},
{-32'd1102, 32'd4926, -32'd1356, 32'd11650},
{32'd10074, -32'd7383, -32'd1364, -32'd1879},
{-32'd2921, 32'd149, 32'd16806, -32'd3139},
{-32'd13119, -32'd14594, -32'd1674, 32'd12546},
{-32'd5014, 32'd8107, 32'd9831, 32'd603},
{-32'd8604, -32'd7640, 32'd3887, -32'd7531},
{32'd1514, 32'd9417, -32'd2508, 32'd12028},
{32'd10174, 32'd284, -32'd9899, 32'd1047},
{-32'd3667, 32'd12558, 32'd624, 32'd7744},
{32'd26224, 32'd10478, 32'd5292, -32'd2416},
{32'd6073, -32'd8642, -32'd3356, 32'd3528},
{32'd1433, -32'd2764, -32'd3643, -32'd2120},
{32'd6855, -32'd1709, -32'd6103, -32'd3160},
{-32'd2611, -32'd10605, 32'd7935, -32'd10336},
{-32'd6863, -32'd1775, -32'd8921, -32'd12299},
{-32'd2527, -32'd3937, -32'd13339, -32'd1409},
{-32'd10552, -32'd15912, 32'd3658, -32'd6044},
{32'd15221, 32'd5199, 32'd6644, 32'd6233},
{32'd897, 32'd14765, 32'd1303, -32'd920},
{-32'd4017, -32'd16199, -32'd8252, 32'd4955},
{-32'd3769, 32'd775, 32'd11799, 32'd4128},
{-32'd4050, 32'd20668, -32'd5310, -32'd4767},
{-32'd11214, -32'd4100, 32'd3913, 32'd1547},
{32'd2956, 32'd1435, -32'd6691, 32'd3622},
{32'd7542, -32'd2657, -32'd3187, -32'd474},
{32'd8702, -32'd13576, -32'd4777, -32'd1506},
{32'd5073, 32'd2623, -32'd8966, -32'd4939},
{32'd473, 32'd680, 32'd18065, 32'd2360},
{-32'd5977, 32'd11956, -32'd8168, 32'd10516},
{-32'd30, -32'd12135, 32'd1696, 32'd1476},
{-32'd8341, -32'd12841, -32'd628, -32'd17181},
{32'd7230, 32'd2132, 32'd6589, -32'd183},
{-32'd8335, 32'd4102, -32'd8627, 32'd5455},
{-32'd6331, 32'd6847, 32'd5817, -32'd2846},
{32'd5858, 32'd12745, 32'd6175, -32'd8395},
{-32'd15438, -32'd4887, 32'd10213, 32'd10706},
{32'd699, 32'd7403, 32'd12286, 32'd4306},
{-32'd4057, -32'd6038, -32'd2922, -32'd6805},
{32'd7190, -32'd13412, 32'd4155, -32'd6703},
{-32'd1542, 32'd5196, -32'd2680, -32'd1828},
{32'd138, -32'd10322, -32'd2000, -32'd5508},
{32'd679, 32'd2454, 32'd5416, 32'd12375},
{32'd8632, 32'd844, -32'd3752, 32'd10347},
{32'd17539, 32'd4619, 32'd8460, -32'd3883},
{32'd7933, -32'd12725, -32'd11483, -32'd22642},
{32'd4838, 32'd7120, -32'd8631, 32'd3062},
{32'd11070, 32'd792, 32'd6331, 32'd6887},
{-32'd3987, 32'd7767, -32'd13308, 32'd3155},
{-32'd6953, 32'd1736, -32'd8142, -32'd4256},
{32'd5883, 32'd2569, 32'd8888, 32'd4440},
{-32'd1250, -32'd9267, 32'd4285, 32'd19136},
{-32'd2479, 32'd6293, -32'd12482, -32'd653},
{-32'd568, 32'd10770, 32'd20383, 32'd1723},
{-32'd957, -32'd9537, 32'd7494, -32'd4192},
{32'd9178, -32'd2526, -32'd4002, 32'd7710},
{32'd924, 32'd11935, -32'd4229, 32'd15964},
{32'd7502, -32'd2833, -32'd3219, -32'd7614},
{32'd1021, 32'd2058, 32'd8039, -32'd2879},
{-32'd14647, -32'd11184, -32'd10868, -32'd5007},
{32'd5237, -32'd3236, -32'd704, 32'd9243},
{-32'd1087, -32'd13116, 32'd5487, -32'd79},
{32'd6194, 32'd509, -32'd4594, -32'd2446},
{32'd3840, 32'd3485, -32'd6219, 32'd10023},
{32'd2473, -32'd6842, -32'd3803, 32'd5419},
{-32'd7333, 32'd7701, 32'd1740, -32'd4632},
{32'd3228, 32'd1037, -32'd5904, -32'd4736},
{32'd2261, -32'd3706, 32'd1329, -32'd9143},
{-32'd13580, -32'd1300, -32'd6369, -32'd1720},
{-32'd5817, 32'd2594, -32'd3356, -32'd1022},
{-32'd5144, 32'd1176, 32'd13399, 32'd14886},
{32'd4432, -32'd6987, 32'd9552, 32'd5664},
{32'd7221, 32'd1503, 32'd3256, -32'd10735},
{32'd12700, -32'd84, -32'd4668, -32'd5411},
{32'd8707, 32'd1233, -32'd6652, 32'd1758},
{32'd5871, 32'd9254, 32'd2421, 32'd2205},
{-32'd7635, -32'd3230, -32'd782, 32'd8277},
{-32'd679, -32'd277, -32'd4464, 32'd9719},
{-32'd10641, -32'd694, 32'd14001, -32'd16991},
{32'd4939, 32'd2113, 32'd1331, 32'd1643},
{32'd835, -32'd10793, -32'd9233, 32'd3989},
{32'd237, 32'd5669, 32'd5799, 32'd13142},
{-32'd14649, -32'd12083, -32'd16016, -32'd699},
{32'd294, 32'd13527, 32'd7235, 32'd15760},
{-32'd1596, 32'd798, -32'd2502, -32'd12411},
{-32'd18475, 32'd11611, -32'd3066, -32'd5869},
{32'd212, 32'd3633, -32'd11401, -32'd1858},
{-32'd10931, -32'd8240, -32'd736, -32'd451},
{32'd8333, 32'd538, -32'd5146, -32'd1077},
{32'd6566, -32'd1091, -32'd7550, 32'd14659},
{32'd10715, 32'd9722, -32'd10601, -32'd5585},
{-32'd1686, 32'd1753, -32'd1185, 32'd15196},
{-32'd10172, -32'd8276, 32'd9085, -32'd2640},
{-32'd8426, -32'd1450, -32'd655, -32'd6999},
{-32'd12949, -32'd7816, 32'd8891, -32'd4310},
{-32'd7030, -32'd13208, -32'd4886, 32'd8155},
{32'd8740, 32'd5832, 32'd1370, -32'd11109},
{32'd13069, -32'd10305, 32'd8946, -32'd683},
{32'd8619, 32'd12223, -32'd1542, 32'd2203},
{32'd9807, 32'd7919, 32'd14664, -32'd12851},
{32'd5168, -32'd1409, -32'd6506, -32'd3932},
{32'd3990, -32'd2669, -32'd6123, 32'd13752},
{32'd139, -32'd7699, 32'd3834, 32'd1534},
{-32'd10560, -32'd2657, -32'd1312, 32'd4288},
{32'd6968, 32'd7560, -32'd11073, 32'd6020},
{32'd13675, 32'd6293, 32'd11571, -32'd2041},
{-32'd4267, 32'd6377, 32'd5210, 32'd843},
{-32'd15906, 32'd2376, 32'd5993, 32'd6190},
{32'd5216, -32'd5406, -32'd15819, -32'd2482},
{-32'd1276, -32'd1647, 32'd5438, 32'd9036},
{-32'd502, -32'd150, 32'd1530, -32'd2754},
{32'd2337, 32'd989, 32'd11255, 32'd4728},
{32'd152, -32'd10993, 32'd3118, -32'd18602},
{-32'd1654, -32'd10392, -32'd9737, 32'd6073},
{32'd2690, 32'd12592, -32'd2769, -32'd4700},
{32'd1914, -32'd5444, 32'd14554, 32'd8275},
{-32'd8745, -32'd22836, 32'd1604, 32'd4124},
{-32'd2097, -32'd1843, 32'd9546, -32'd5994},
{-32'd6191, 32'd2664, -32'd7587, -32'd6762},
{-32'd14187, -32'd5648, 32'd1229, -32'd10248},
{-32'd1418, -32'd3921, 32'd6028, -32'd433},
{-32'd2643, 32'd4848, -32'd9282, 32'd824},
{-32'd2376, 32'd5616, -32'd2100, -32'd12872},
{32'd8628, -32'd1316, -32'd12576, 32'd1637},
{32'd1762, -32'd6172, -32'd16048, -32'd10600},
{-32'd9679, -32'd2089, 32'd1535, 32'd19300},
{-32'd1595, 32'd4739, -32'd433, -32'd2401},
{32'd8797, -32'd9727, -32'd3590, -32'd3066},
{-32'd9599, 32'd2444, 32'd2350, 32'd4029},
{32'd14828, 32'd2199, -32'd12784, -32'd2418},
{-32'd8365, 32'd17006, -32'd3951, -32'd8799},
{32'd5002, -32'd7747, 32'd3246, 32'd1649},
{32'd11329, -32'd4022, 32'd2911, 32'd1137},
{-32'd5687, 32'd400, 32'd1951, 32'd5570},
{32'd5549, 32'd4867, -32'd338, -32'd613},
{-32'd1156, -32'd2200, -32'd3397, -32'd9528},
{-32'd4944, -32'd10210, -32'd3628, -32'd19564},
{32'd4053, 32'd13806, -32'd5248, -32'd1433},
{32'd2840, 32'd4367, 32'd4719, 32'd6547},
{32'd10261, -32'd7850, -32'd1736, -32'd5715},
{-32'd2757, 32'd216, 32'd12919, 32'd3812},
{32'd11164, -32'd10960, 32'd89, -32'd4587},
{32'd6703, -32'd1434, 32'd3896, -32'd10666},
{32'd7833, -32'd2004, -32'd1121, 32'd5852},
{32'd9977, -32'd7418, 32'd1521, 32'd4879},
{-32'd2489, -32'd5166, -32'd6612, -32'd5719},
{32'd7713, -32'd4919, -32'd3719, -32'd6614},
{32'd6582, -32'd5424, 32'd3067, 32'd14008},
{-32'd5768, -32'd977, -32'd980, 32'd9227},
{-32'd3856, 32'd2226, 32'd9074, 32'd1075},
{-32'd3334, -32'd4415, 32'd3048, -32'd1508},
{-32'd6603, -32'd874, -32'd8870, -32'd5971},
{32'd10388, 32'd25290, 32'd3346, 32'd9227},
{32'd14515, 32'd9832, -32'd4089, 32'd2464},
{32'd4252, 32'd2897, -32'd12423, 32'd417},
{32'd4689, 32'd5769, 32'd15494, -32'd5049},
{32'd683, 32'd2049, 32'd4418, -32'd2699},
{32'd7780, 32'd1005, 32'd15247, -32'd212},
{-32'd7931, -32'd11340, -32'd2273, -32'd10326},
{-32'd8844, -32'd352, 32'd6545, 32'd4465},
{-32'd12903, 32'd13781, 32'd9770, 32'd5727},
{32'd6171, -32'd3766, -32'd8021, -32'd1006},
{32'd5466, 32'd12090, 32'd1507, 32'd1027},
{32'd7338, 32'd141, 32'd4163, 32'd8209},
{32'd10628, -32'd3087, -32'd12939, -32'd2306},
{32'd6693, -32'd8282, 32'd7681, -32'd50},
{-32'd7110, -32'd9326, -32'd3154, 32'd3008},
{-32'd8919, 32'd7876, 32'd6256, -32'd4720},
{-32'd8177, -32'd683, -32'd6485, -32'd2930},
{32'd12445, -32'd19229, 32'd5088, 32'd1856},
{-32'd3906, 32'd3688, -32'd5225, -32'd6716},
{-32'd9012, -32'd9957, 32'd6393, -32'd1372},
{-32'd7126, -32'd3695, 32'd7798, 32'd5066},
{-32'd431, 32'd2549, -32'd4676, -32'd3322},
{32'd13128, -32'd988, -32'd5121, -32'd8535},
{32'd11688, -32'd9184, 32'd14651, -32'd3419},
{-32'd9844, -32'd13589, -32'd4054, 32'd1205},
{-32'd5607, -32'd5278, 32'd6088, -32'd2294},
{32'd1662, 32'd10414, -32'd3431, -32'd1356},
{32'd5550, 32'd8530, -32'd6660, -32'd6928},
{32'd2173, 32'd4917, 32'd11104, -32'd4596},
{-32'd7174, -32'd14405, -32'd4551, 32'd2443},
{32'd1253, 32'd5240, -32'd3780, 32'd6562},
{32'd1795, 32'd1833, 32'd4568, -32'd1049},
{32'd4507, 32'd1484, 32'd1024, -32'd4505},
{-32'd14203, 32'd64, -32'd1299, -32'd4929},
{-32'd6304, -32'd1323, 32'd590, -32'd2724},
{32'd14561, -32'd4934, 32'd3383, 32'd6276},
{32'd9540, -32'd1770, -32'd6351, 32'd3721},
{32'd9983, 32'd2330, -32'd10615, -32'd6120},
{-32'd623, -32'd1471, -32'd559, -32'd2615},
{-32'd3553, 32'd2373, -32'd3327, -32'd14772},
{-32'd14066, 32'd3921, 32'd3513, 32'd4671},
{32'd7558, -32'd2110, -32'd12212, -32'd4814},
{32'd4960, 32'd4797, -32'd17072, 32'd205},
{-32'd246, -32'd2528, -32'd586, 32'd13886},
{-32'd5017, -32'd5149, -32'd19399, 32'd7735},
{-32'd3573, -32'd6715, -32'd3205, 32'd6645},
{32'd2931, 32'd10384, 32'd12389, 32'd5461},
{-32'd7561, 32'd10468, -32'd7669, -32'd8193},
{32'd1502, -32'd8785, -32'd7113, 32'd9327},
{32'd5615, -32'd7384, 32'd15354, 32'd11731},
{-32'd1107, 32'd4045, -32'd5950, -32'd2925},
{32'd3008, -32'd9261, -32'd1300, -32'd6623},
{-32'd5838, 32'd9217, 32'd2213, -32'd17067},
{32'd7106, -32'd4233, -32'd7313, -32'd7510},
{32'd6232, -32'd1944, 32'd6060, 32'd18437},
{-32'd795, 32'd1468, 32'd8707, -32'd6892},
{-32'd3980, 32'd1578, 32'd4278, -32'd9726},
{32'd3476, 32'd1283, -32'd2504, -32'd1368},
{-32'd6123, -32'd708, -32'd2139, -32'd11819},
{32'd3693, -32'd11879, -32'd10688, 32'd6763},
{32'd12311, 32'd161, -32'd17139, -32'd3656},
{-32'd682, -32'd2318, -32'd11797, -32'd2532},
{32'd18266, -32'd3251, 32'd6168, 32'd4510},
{32'd3753, 32'd118, -32'd7237, 32'd2224},
{-32'd5533, -32'd3592, -32'd1364, -32'd3597},
{-32'd10541, 32'd12990, -32'd7178, -32'd3367},
{32'd1020, 32'd10779, 32'd8052, -32'd454},
{-32'd266, 32'd3997, -32'd4816, -32'd4368},
{-32'd10585, -32'd2046, -32'd2681, 32'd2436},
{32'd14294, -32'd5210, -32'd6613, -32'd471},
{32'd14675, 32'd3516, 32'd779, -32'd5753},
{32'd4218, -32'd5698, 32'd3655, 32'd3653},
{-32'd6514, -32'd7671, -32'd2152, -32'd6726},
{-32'd2007, -32'd2288, 32'd7415, 32'd4159},
{-32'd513, 32'd1402, 32'd5853, -32'd8261},
{-32'd4384, -32'd1346, 32'd6860, 32'd17527},
{32'd15192, 32'd11313, 32'd12523, -32'd9401},
{-32'd11347, -32'd18422, -32'd6772, -32'd4355},
{32'd1730, 32'd5596, 32'd9060, 32'd2807},
{-32'd15587, -32'd248, -32'd670, -32'd6691},
{-32'd3985, -32'd3438, -32'd14575, -32'd400},
{32'd4348, -32'd1004, -32'd11436, 32'd2153},
{32'd12808, 32'd2110, -32'd3448, 32'd18149},
{-32'd11579, 32'd2561, 32'd5733, -32'd785},
{32'd3613, 32'd6979, -32'd2234, -32'd5533},
{-32'd12956, 32'd3937, -32'd8607, -32'd10241},
{32'd2561, 32'd12490, -32'd5874, 32'd8599},
{32'd3951, -32'd818, -32'd7768, 32'd10003},
{-32'd5403, -32'd933, 32'd11526, 32'd10713},
{32'd5277, -32'd12264, -32'd16087, -32'd11244},
{32'd11238, 32'd1411, -32'd9531, -32'd6544},
{32'd5730, -32'd13939, 32'd2576, 32'd10642},
{-32'd13172, -32'd9323, -32'd3598, 32'd605},
{-32'd1006, 32'd13055, 32'd12793, -32'd1611},
{-32'd12049, -32'd8431, 32'd6315, 32'd3635},
{-32'd2913, -32'd7483, 32'd8134, -32'd15991},
{-32'd1116, -32'd2650, -32'd13748, -32'd3348},
{32'd8494, -32'd3592, -32'd15963, 32'd4588},
{32'd11883, 32'd5137, -32'd2282, -32'd14762},
{32'd2169, 32'd6823, -32'd770, 32'd1656},
{-32'd5467, -32'd1875, -32'd2182, -32'd194},
{32'd2206, -32'd2391, 32'd1930, -32'd11963}
},
{{32'd15363, 32'd12888, 32'd8401, -32'd2277},
{32'd1619, -32'd15745, -32'd2507, 32'd102},
{32'd800, 32'd6322, 32'd403, -32'd3117},
{32'd1735, -32'd1452, 32'd4765, 32'd9952},
{-32'd6115, -32'd11066, -32'd7378, 32'd3968},
{-32'd10874, 32'd841, 32'd6868, -32'd2167},
{32'd5999, 32'd9161, 32'd1169, 32'd1602},
{-32'd1574, -32'd15798, 32'd4261, -32'd6132},
{32'd7129, 32'd9172, -32'd4077, 32'd10376},
{32'd8410, 32'd2479, 32'd9795, 32'd4997},
{-32'd877, 32'd6204, -32'd6281, -32'd5755},
{32'd4756, -32'd7606, 32'd1422, -32'd9017},
{32'd129, 32'd904, -32'd694, 32'd6735},
{-32'd6216, -32'd12425, -32'd7492, 32'd6858},
{32'd1199, -32'd2813, -32'd3586, 32'd7657},
{32'd7668, 32'd1788, -32'd9332, 32'd1842},
{-32'd3044, -32'd1092, 32'd3840, 32'd1948},
{-32'd4245, -32'd6795, 32'd3288, 32'd228},
{32'd5226, -32'd3624, 32'd255, 32'd4339},
{32'd5259, 32'd14935, -32'd1861, 32'd7812},
{-32'd4181, -32'd2572, -32'd8233, 32'd1360},
{-32'd14676, 32'd1521, 32'd2822, 32'd13272},
{-32'd8367, -32'd9084, -32'd5803, -32'd223},
{-32'd9832, 32'd1654, 32'd8340, -32'd5650},
{32'd4455, 32'd14683, 32'd1772, -32'd4170},
{-32'd4283, 32'd7281, 32'd7117, -32'd4028},
{-32'd6821, 32'd12063, -32'd1323, -32'd4047},
{32'd3838, -32'd2394, 32'd3572, 32'd1332},
{-32'd263, -32'd10508, 32'd9974, -32'd7506},
{32'd514, 32'd4498, -32'd16580, 32'd958},
{32'd410, 32'd11590, 32'd4975, 32'd14494},
{-32'd6374, -32'd5128, 32'd1126, -32'd396},
{32'd2624, -32'd5689, -32'd1591, -32'd5154},
{-32'd12688, 32'd2417, -32'd9270, -32'd901},
{-32'd2433, 32'd3934, 32'd6813, 32'd8028},
{32'd8976, 32'd9995, 32'd4926, -32'd5906},
{-32'd7293, -32'd2653, -32'd5775, 32'd5502},
{32'd6572, -32'd749, -32'd861, 32'd1723},
{-32'd6469, -32'd7334, -32'd164, 32'd7827},
{32'd1055, 32'd13678, 32'd13103, -32'd3583},
{-32'd3305, -32'd1296, 32'd231, -32'd7519},
{-32'd1459, 32'd13548, -32'd380, 32'd2157},
{32'd7656, -32'd8063, 32'd1069, 32'd6183},
{-32'd1092, -32'd12144, -32'd2194, 32'd437},
{-32'd8397, 32'd4102, 32'd6352, 32'd7995},
{32'd10469, -32'd5582, -32'd2256, 32'd1320},
{32'd807, -32'd3928, 32'd2294, 32'd263},
{-32'd6755, -32'd12211, -32'd10401, -32'd4163},
{32'd15766, 32'd7804, -32'd12721, 32'd9222},
{32'd8783, -32'd8130, 32'd5869, 32'd2835},
{-32'd9392, 32'd3317, 32'd9760, -32'd1349},
{32'd6275, 32'd1344, -32'd5124, -32'd2001},
{-32'd15223, -32'd13110, -32'd4578, 32'd7791},
{32'd3080, -32'd9863, 32'd2464, 32'd3813},
{32'd2858, -32'd2310, 32'd4908, 32'd2200},
{-32'd7992, 32'd2285, 32'd3084, -32'd8435},
{32'd11768, 32'd5456, 32'd9555, 32'd2845},
{-32'd10569, 32'd894, -32'd4421, 32'd1937},
{32'd14831, -32'd9085, 32'd6250, -32'd1617},
{32'd293, 32'd5840, -32'd10731, -32'd10579},
{-32'd21348, -32'd2207, 32'd8312, 32'd6962},
{32'd6962, 32'd2245, 32'd6967, 32'd2217},
{32'd943, -32'd462, 32'd3749, 32'd70},
{-32'd49, -32'd1821, -32'd1143, 32'd309},
{-32'd8039, -32'd11, -32'd3594, 32'd869},
{32'd3654, 32'd14517, 32'd10077, 32'd7150},
{-32'd7503, -32'd9682, -32'd1226, -32'd6401},
{32'd488, -32'd3089, -32'd2761, 32'd6748},
{32'd7239, -32'd386, -32'd2893, -32'd8972},
{-32'd7759, 32'd10069, 32'd6541, -32'd6207},
{32'd2007, -32'd14719, -32'd7669, -32'd2607},
{-32'd6518, 32'd5099, -32'd1856, 32'd1186},
{-32'd15179, 32'd8493, 32'd1165, 32'd258},
{32'd1842, 32'd2624, -32'd8662, -32'd635},
{-32'd13594, 32'd7856, 32'd831, -32'd4157},
{32'd10683, -32'd2394, 32'd1684, 32'd1088},
{-32'd2995, -32'd17481, -32'd12345, -32'd5308},
{32'd4329, 32'd5922, -32'd8006, -32'd7625},
{32'd207, -32'd1775, -32'd1826, 32'd7930},
{32'd40, -32'd10393, 32'd9022, -32'd2108},
{32'd8318, 32'd1343, -32'd12671, -32'd13785},
{32'd1055, 32'd696, -32'd4574, 32'd8197},
{-32'd10825, -32'd9786, -32'd118, -32'd68},
{-32'd4769, -32'd4873, -32'd3630, -32'd5588},
{32'd1132, -32'd10382, -32'd1370, -32'd1106},
{-32'd9994, 32'd3891, 32'd11088, -32'd3556},
{-32'd2518, 32'd7151, -32'd3815, -32'd2790},
{-32'd3936, -32'd4154, -32'd6261, 32'd4329},
{32'd14370, -32'd7789, -32'd4666, 32'd2846},
{32'd3716, -32'd13929, -32'd11448, -32'd2891},
{32'd17378, 32'd3375, 32'd6336, 32'd5919},
{-32'd2275, 32'd12649, -32'd435, -32'd87},
{32'd2582, -32'd5487, -32'd579, 32'd6519},
{-32'd7699, -32'd11433, -32'd9415, 32'd6414},
{-32'd7109, -32'd473, 32'd10368, -32'd2461},
{-32'd2762, -32'd2326, -32'd9179, 32'd1048},
{32'd4165, -32'd7026, 32'd6585, 32'd5944},
{-32'd6296, -32'd5813, 32'd6301, -32'd173},
{32'd364, 32'd3292, 32'd4957, 32'd3946},
{32'd6493, -32'd3864, -32'd6146, 32'd8597},
{-32'd3334, -32'd6671, -32'd9293, -32'd3184},
{32'd2259, 32'd5727, 32'd2302, -32'd7484},
{32'd7978, -32'd1344, 32'd480, 32'd3080},
{32'd13901, -32'd8577, 32'd538, -32'd6224},
{32'd2953, 32'd4200, 32'd5755, 32'd5975},
{32'd1591, 32'd4898, -32'd3729, -32'd9762},
{32'd2333, -32'd2318, -32'd5676, -32'd5980},
{-32'd4510, -32'd13221, 32'd863, -32'd1401},
{32'd851, -32'd3189, 32'd1008, 32'd264},
{32'd9358, 32'd1364, 32'd7141, -32'd754},
{-32'd4767, -32'd7902, -32'd13451, -32'd1848},
{-32'd11972, 32'd3169, -32'd5166, -32'd3988},
{-32'd3687, 32'd986, 32'd7853, 32'd7499},
{-32'd17890, 32'd6310, 32'd449, -32'd1676},
{-32'd3672, -32'd7915, -32'd14645, -32'd9562},
{32'd7117, 32'd11713, -32'd11196, 32'd97},
{-32'd6170, 32'd981, 32'd3804, -32'd1080},
{32'd7273, 32'd91, -32'd152, -32'd8115},
{-32'd3859, -32'd1738, 32'd5726, -32'd6862},
{32'd320, 32'd912, 32'd6606, 32'd18320},
{32'd7450, 32'd1474, 32'd4550, 32'd9922},
{-32'd11299, 32'd3055, 32'd4141, 32'd8338},
{32'd5894, -32'd13141, -32'd3974, 32'd4135},
{-32'd750, -32'd1741, 32'd780, -32'd12885},
{-32'd17406, 32'd3329, -32'd8244, 32'd7702},
{-32'd5883, -32'd4684, 32'd18928, 32'd3511},
{-32'd6424, 32'd6971, -32'd2821, 32'd3438},
{-32'd6250, -32'd16669, 32'd4737, 32'd8476},
{-32'd3803, 32'd3463, -32'd3719, -32'd6976},
{-32'd2147, 32'd3031, 32'd7592, 32'd3166},
{32'd1219, 32'd8279, 32'd3286, 32'd5084},
{32'd5682, -32'd9818, 32'd5842, -32'd5477},
{-32'd8619, 32'd1311, -32'd6741, 32'd396},
{32'd8631, -32'd8204, 32'd8596, -32'd5231},
{-32'd10659, 32'd3884, 32'd4057, 32'd2573},
{-32'd3994, -32'd1439, 32'd4475, -32'd5661},
{32'd1309, 32'd2204, -32'd566, 32'd2603},
{32'd6740, -32'd10549, -32'd6022, -32'd1854},
{32'd5659, -32'd7044, -32'd4806, -32'd4511},
{32'd4747, -32'd6395, -32'd11110, -32'd12904},
{-32'd4150, 32'd10960, -32'd8420, 32'd149},
{32'd9384, -32'd7542, -32'd452, -32'd693},
{32'd6745, 32'd625, 32'd1849, 32'd8241},
{32'd7748, 32'd6816, 32'd2050, -32'd694},
{-32'd7305, 32'd6438, -32'd5752, 32'd3638},
{32'd8091, -32'd2312, -32'd13604, 32'd3627},
{-32'd8706, -32'd843, 32'd9245, 32'd9401},
{32'd3153, 32'd6492, 32'd9924, 32'd3596},
{32'd3389, 32'd7293, 32'd1332, 32'd4753},
{-32'd625, -32'd5280, -32'd930, 32'd1986},
{32'd7396, -32'd1126, -32'd15165, 32'd529},
{-32'd5212, -32'd10398, 32'd5788, 32'd7332},
{32'd4160, -32'd4650, -32'd8481, 32'd5382},
{-32'd13517, -32'd3751, -32'd9072, 32'd2369},
{32'd2026, 32'd2428, -32'd2843, -32'd4979},
{-32'd7798, -32'd15615, -32'd9519, 32'd5020},
{32'd5189, 32'd11145, 32'd8085, 32'd11237},
{-32'd15288, -32'd1234, 32'd15655, 32'd3615},
{-32'd13716, -32'd10850, -32'd3029, 32'd2839},
{32'd14150, 32'd14140, -32'd2422, 32'd3581},
{32'd3003, -32'd6315, -32'd2620, 32'd1111},
{-32'd1967, 32'd3180, 32'd10637, 32'd32},
{-32'd12638, 32'd4629, -32'd8074, -32'd3567},
{-32'd2943, -32'd2847, 32'd14849, 32'd2945},
{32'd16164, 32'd5477, -32'd4950, 32'd1875},
{-32'd2560, -32'd8011, -32'd3110, -32'd10097},
{32'd9431, 32'd3990, -32'd1587, 32'd4829},
{-32'd3635, -32'd2886, 32'd12215, -32'd583},
{-32'd11866, 32'd3285, -32'd2248, -32'd6457},
{-32'd8920, 32'd4237, -32'd6691, 32'd2596},
{32'd2956, -32'd1712, -32'd2058, -32'd4437},
{32'd4319, -32'd2355, -32'd14266, -32'd4971},
{32'd3213, 32'd4650, 32'd8712, -32'd6146},
{32'd870, 32'd1163, -32'd2419, -32'd339},
{32'd4859, 32'd166, 32'd2683, 32'd524},
{-32'd1248, 32'd2219, 32'd5252, 32'd2539},
{-32'd2212, -32'd10519, 32'd6920, -32'd4917},
{-32'd3070, -32'd139, -32'd619, -32'd2122},
{32'd21505, -32'd628, 32'd12502, 32'd3876},
{32'd3060, -32'd11171, -32'd6158, -32'd3164},
{-32'd841, -32'd6361, -32'd12709, -32'd2737},
{32'd8454, -32'd9232, -32'd7225, 32'd15351},
{32'd15493, 32'd1688, -32'd8640, -32'd2201},
{32'd7999, 32'd9788, -32'd17726, 32'd6961},
{32'd6124, -32'd6635, 32'd659, 32'd1087},
{-32'd9048, 32'd2455, -32'd1717, -32'd83},
{32'd1219, 32'd7088, 32'd11589, -32'd1393},
{32'd4068, -32'd5864, -32'd1822, 32'd1377},
{-32'd235, -32'd4499, 32'd2914, 32'd6838},
{-32'd10184, -32'd14457, 32'd1924, -32'd6826},
{-32'd7158, -32'd102, 32'd6709, 32'd8661},
{32'd10574, -32'd7514, -32'd1565, 32'd2234},
{32'd3184, -32'd8261, -32'd2655, -32'd4795},
{32'd3823, 32'd7085, 32'd4391, 32'd9355},
{-32'd4593, -32'd3228, -32'd4896, 32'd3347},
{-32'd4568, 32'd3686, -32'd10138, -32'd7247},
{32'd2398, 32'd1547, -32'd5209, -32'd14115},
{32'd4952, 32'd18211, 32'd5727, 32'd3750},
{-32'd3133, -32'd6785, 32'd8143, -32'd6254},
{32'd7259, -32'd2404, -32'd71, -32'd530},
{32'd3240, -32'd3029, -32'd9300, -32'd3738},
{-32'd6285, 32'd10188, -32'd9140, -32'd5838},
{32'd5486, 32'd1089, -32'd1461, 32'd3803},
{-32'd6270, -32'd5624, -32'd55, -32'd2554},
{-32'd11132, -32'd2260, 32'd3146, 32'd566},
{32'd2918, -32'd5579, 32'd950, -32'd5089},
{32'd6334, 32'd1792, -32'd10653, 32'd3250},
{32'd3207, -32'd4725, -32'd18933, 32'd1397},
{-32'd8286, 32'd2520, 32'd919, -32'd1221},
{32'd17960, -32'd5672, -32'd4431, 32'd3252},
{-32'd3562, 32'd10120, -32'd16031, -32'd3560},
{32'd7320, 32'd1793, -32'd13696, 32'd9171},
{-32'd10986, 32'd6062, 32'd9689, -32'd5930},
{32'd4582, -32'd96, -32'd10751, -32'd457},
{32'd3638, 32'd13063, -32'd4363, 32'd5054},
{-32'd12711, -32'd203, -32'd1820, -32'd2075},
{-32'd6661, 32'd1921, -32'd859, -32'd6556},
{-32'd4553, -32'd2281, -32'd4040, -32'd2919},
{32'd5268, 32'd3775, 32'd5655, -32'd1110},
{-32'd9954, 32'd11457, 32'd5143, -32'd8803},
{32'd13895, -32'd4210, -32'd8348, 32'd3122},
{-32'd8928, 32'd8020, 32'd6446, -32'd3503},
{32'd3735, 32'd1857, 32'd3739, 32'd4513},
{32'd2372, 32'd3368, -32'd3602, -32'd12021},
{32'd6270, -32'd6216, 32'd399, -32'd5135},
{32'd13521, -32'd1154, 32'd3069, 32'd291},
{32'd3627, 32'd2993, 32'd8124, -32'd2270},
{32'd1246, 32'd1540, 32'd7846, -32'd4612},
{32'd8235, 32'd7528, -32'd14317, 32'd2540},
{-32'd8931, 32'd1871, 32'd12031, 32'd8589},
{32'd1945, 32'd8870, -32'd12285, -32'd5399},
{-32'd3904, 32'd5550, -32'd7849, -32'd11185},
{32'd7158, 32'd8509, 32'd3750, -32'd5048},
{-32'd10188, -32'd920, -32'd7399, -32'd5490},
{32'd4105, -32'd12120, 32'd6735, -32'd5062},
{-32'd4201, -32'd327, -32'd11272, 32'd3165},
{32'd6882, -32'd6256, -32'd7884, 32'd4568},
{-32'd9805, 32'd679, 32'd7963, -32'd1821},
{32'd14802, -32'd2442, 32'd6814, -32'd8717},
{32'd4174, -32'd3626, -32'd3829, 32'd3489},
{-32'd8955, 32'd14167, 32'd4222, -32'd4796},
{-32'd804, 32'd8811, -32'd5110, -32'd5767},
{32'd288, -32'd10232, -32'd5283, -32'd1570},
{-32'd10696, 32'd12739, 32'd4360, 32'd2369},
{32'd419, 32'd2962, -32'd799, -32'd2464},
{-32'd14871, -32'd3460, -32'd12046, -32'd5874},
{32'd351, -32'd9261, -32'd1086, -32'd5934},
{-32'd10596, -32'd8517, 32'd4008, -32'd11677},
{32'd849, -32'd13787, -32'd5133, -32'd6562},
{32'd5454, -32'd1945, 32'd11583, -32'd2153},
{-32'd6436, 32'd4215, -32'd6815, -32'd6270},
{-32'd3960, -32'd1300, -32'd2958, -32'd6102},
{-32'd13494, -32'd698, -32'd2773, -32'd5622},
{-32'd2829, -32'd6635, -32'd2516, 32'd4059},
{-32'd2423, 32'd1031, -32'd9614, 32'd3452},
{-32'd8974, -32'd2543, -32'd2829, -32'd3187},
{32'd776, 32'd227, -32'd9906, 32'd4991},
{32'd2534, 32'd1961, 32'd4897, 32'd13909},
{32'd2329, -32'd2416, -32'd2252, -32'd1904},
{32'd3514, -32'd1881, -32'd2925, -32'd3721},
{-32'd13387, 32'd875, 32'd400, -32'd6860},
{-32'd11342, -32'd7390, -32'd2595, -32'd4591},
{-32'd9972, 32'd2795, -32'd17697, -32'd3430},
{-32'd1467, 32'd9378, -32'd6345, -32'd13098},
{-32'd2351, 32'd9397, -32'd4270, 32'd7051},
{-32'd6267, -32'd4442, 32'd13033, -32'd1627},
{32'd4952, -32'd2272, 32'd3422, 32'd1637},
{-32'd11114, 32'd15426, 32'd11165, 32'd14569},
{-32'd7932, -32'd7045, -32'd7, 32'd5379},
{-32'd4019, 32'd3444, -32'd5998, -32'd5764},
{32'd7877, -32'd5202, -32'd5121, -32'd5572},
{-32'd1304, 32'd8815, -32'd1018, 32'd622},
{-32'd6974, -32'd15060, 32'd691, 32'd771},
{32'd9040, -32'd3596, -32'd2727, -32'd3781},
{32'd10783, -32'd14533, 32'd180, -32'd504},
{-32'd7483, 32'd1603, 32'd3235, 32'd264},
{32'd2349, 32'd3408, 32'd10410, 32'd5983},
{32'd5153, 32'd16326, -32'd590, -32'd86},
{-32'd5810, -32'd3499, 32'd6356, -32'd5259},
{-32'd1633, -32'd7975, 32'd11849, 32'd8460},
{-32'd10614, -32'd1107, 32'd12722, 32'd554},
{32'd9021, 32'd3161, 32'd211, 32'd1082},
{32'd14503, 32'd342, -32'd6348, -32'd975},
{32'd6242, -32'd495, 32'd10725, -32'd6204},
{32'd2532, 32'd2380, 32'd1991, 32'd1698},
{-32'd2511, -32'd9409, -32'd1689, -32'd2083},
{-32'd4389, -32'd5960, -32'd1000, 32'd2894},
{-32'd14551, 32'd8875, -32'd6248, 32'd1690},
{32'd3933, -32'd1827, -32'd2069, -32'd1661},
{-32'd13995, -32'd7869, 32'd4188, -32'd236},
{-32'd4276, 32'd3762, 32'd657, 32'd13541},
{32'd11526, -32'd739, -32'd120, 32'd4384},
{-32'd3034, 32'd6271, 32'd4823, -32'd2299},
{-32'd5439, -32'd1545, -32'd1584, -32'd7168},
{32'd7753, -32'd6820, 32'd7635, -32'd9130},
{32'd8078, -32'd4235, -32'd5686, 32'd109},
{-32'd5828, -32'd737, -32'd119, 32'd8524},
{-32'd10623, 32'd7525, -32'd2975, -32'd1131},
{32'd3904, -32'd4399, 32'd299, 32'd910},
{32'd4133, -32'd1030, -32'd2073, 32'd6652}
},
{{-32'd14986, 32'd5555, 32'd6365, 32'd12366},
{32'd8762, -32'd11653, 32'd4507, -32'd9258},
{32'd9855, -32'd10457, 32'd3679, 32'd11096},
{32'd2786, -32'd1001, -32'd6952, 32'd11441},
{32'd8780, -32'd7314, 32'd19789, 32'd23859},
{-32'd687, -32'd212, -32'd10521, 32'd1462},
{-32'd3986, -32'd1941, -32'd742, 32'd9510},
{-32'd3955, 32'd4546, -32'd11783, 32'd6556},
{32'd2924, -32'd10119, 32'd4946, -32'd6592},
{32'd6256, 32'd2848, 32'd3109, 32'd4529},
{32'd8618, -32'd5881, -32'd4082, -32'd8519},
{-32'd4575, -32'd3548, 32'd7184, 32'd5760},
{32'd12436, 32'd1003, 32'd10862, 32'd1165},
{-32'd9724, 32'd7472, -32'd5459, 32'd1327},
{-32'd6034, -32'd3911, 32'd1260, -32'd7121},
{-32'd11898, 32'd11126, 32'd6339, -32'd5663},
{-32'd2549, 32'd11524, 32'd12449, 32'd9546},
{-32'd13985, 32'd3461, -32'd10521, -32'd3647},
{32'd12281, -32'd13947, 32'd325, 32'd4862},
{32'd14791, -32'd8275, 32'd7161, 32'd6220},
{32'd3629, -32'd6386, 32'd4401, -32'd9321},
{32'd2367, -32'd9932, 32'd708, -32'd456},
{-32'd3297, -32'd1984, -32'd7616, 32'd6788},
{-32'd10690, 32'd433, -32'd2523, -32'd10576},
{-32'd915, -32'd3532, 32'd1524, 32'd1312},
{-32'd11211, 32'd11687, -32'd6600, -32'd3355},
{32'd663, -32'd10653, -32'd4141, 32'd180},
{32'd6140, -32'd1368, 32'd2510, -32'd4029},
{-32'd1109, 32'd22430, 32'd4068, 32'd3733},
{-32'd1053, 32'd613, 32'd10319, 32'd808},
{32'd8051, -32'd5264, 32'd729, 32'd1163},
{-32'd3136, -32'd4833, -32'd5184, 32'd3048},
{32'd6132, 32'd18969, -32'd1667, 32'd1998},
{-32'd10103, 32'd1693, 32'd3564, -32'd2518},
{32'd3946, 32'd7449, 32'd11377, 32'd5626},
{-32'd7227, -32'd13521, -32'd360, -32'd954},
{-32'd5806, 32'd1490, 32'd2052, -32'd2757},
{-32'd16880, 32'd17099, -32'd4581, 32'd1302},
{32'd304, 32'd1845, -32'd2354, 32'd5377},
{32'd2877, -32'd1717, -32'd1704, 32'd10918},
{32'd9310, -32'd11597, -32'd5382, -32'd9211},
{-32'd6389, -32'd3141, 32'd6397, -32'd4536},
{-32'd4972, 32'd6594, 32'd1862, 32'd13356},
{-32'd5535, 32'd1424, 32'd4386, -32'd4012},
{-32'd1866, -32'd8527, 32'd888, -32'd4347},
{-32'd3373, -32'd1005, 32'd7504, -32'd4997},
{32'd8511, -32'd14910, -32'd12618, -32'd13233},
{-32'd2761, 32'd2762, -32'd5133, 32'd904},
{-32'd2216, -32'd4378, -32'd1580, -32'd2794},
{-32'd5484, -32'd9161, -32'd4982, 32'd10777},
{-32'd4282, -32'd21138, 32'd9262, 32'd11531},
{-32'd5758, 32'd2022, -32'd1392, -32'd7523},
{-32'd4221, -32'd7856, -32'd9591, 32'd5436},
{32'd9099, 32'd2284, 32'd2499, 32'd3221},
{-32'd3596, 32'd8663, 32'd7380, 32'd5572},
{-32'd5106, -32'd3728, 32'd5084, 32'd2219},
{32'd3103, -32'd4179, -32'd11749, 32'd12899},
{-32'd11911, -32'd759, 32'd1410, -32'd2591},
{32'd5731, -32'd4070, -32'd4291, -32'd4558},
{-32'd5241, -32'd7777, -32'd12840, 32'd10966},
{32'd6593, -32'd17169, 32'd721, 32'd20703},
{32'd262, 32'd3800, 32'd3549, -32'd8066},
{32'd8075, -32'd4669, 32'd8667, -32'd12556},
{32'd4672, -32'd6750, -32'd3444, -32'd2800},
{-32'd6684, -32'd10963, 32'd2709, -32'd13483},
{32'd2769, -32'd6970, -32'd3795, 32'd14038},
{-32'd16598, 32'd10673, 32'd1562, -32'd1642},
{32'd6548, -32'd13536, 32'd8635, -32'd11200},
{-32'd5042, -32'd11514, 32'd2332, -32'd8268},
{-32'd8448, 32'd3668, 32'd5559, -32'd11060},
{-32'd3597, -32'd10128, 32'd809, -32'd4689},
{32'd2396, -32'd1927, 32'd5630, 32'd480},
{-32'd7595, -32'd8421, -32'd13555, -32'd12158},
{32'd2568, -32'd11315, 32'd7383, -32'd5105},
{32'd7445, 32'd11534, 32'd70, 32'd5345},
{-32'd92, -32'd2397, 32'd5646, -32'd1450},
{32'd8917, 32'd11655, -32'd4601, -32'd5144},
{-32'd19395, 32'd7608, 32'd5424, 32'd3090},
{32'd4169, 32'd20865, -32'd4244, -32'd3164},
{32'd1205, 32'd13956, 32'd5816, 32'd855},
{-32'd3371, 32'd10422, -32'd5664, 32'd4110},
{32'd4358, -32'd10877, -32'd1775, 32'd11222},
{32'd12367, 32'd3213, 32'd1037, 32'd3525},
{32'd3706, 32'd9565, 32'd4061, 32'd7983},
{-32'd2694, -32'd2661, 32'd5317, 32'd8373},
{32'd1802, -32'd22274, 32'd413, -32'd17030},
{32'd6586, -32'd5997, 32'd9791, 32'd9829},
{-32'd6845, -32'd8567, 32'd52, -32'd20818},
{32'd3797, 32'd8556, -32'd10193, -32'd11111},
{-32'd434, -32'd1106, -32'd13592, 32'd3333},
{32'd411, -32'd4203, -32'd7872, 32'd8026},
{-32'd8922, -32'd24607, -32'd4409, -32'd1833},
{-32'd3573, 32'd2736, -32'd9108, -32'd8217},
{32'd6759, 32'd20096, 32'd2867, 32'd1223},
{32'd6908, 32'd6607, -32'd3940, -32'd6066},
{32'd4562, -32'd1142, 32'd283, -32'd950},
{-32'd3756, 32'd6351, 32'd7853, 32'd7668},
{-32'd2427, -32'd5841, -32'd13414, 32'd1276},
{-32'd11495, 32'd4796, -32'd2454, -32'd5593},
{-32'd1635, 32'd3286, -32'd6611, 32'd10368},
{32'd16735, -32'd2564, -32'd15612, -32'd17668},
{32'd4910, -32'd14395, 32'd3866, -32'd6823},
{32'd16667, 32'd5326, 32'd3939, -32'd2126},
{-32'd6564, 32'd5776, 32'd10540, -32'd330},
{-32'd895, 32'd18136, -32'd6025, 32'd4687},
{32'd4497, 32'd1503, -32'd4347, -32'd6258},
{32'd6255, -32'd1901, -32'd7903, 32'd1790},
{-32'd8128, 32'd6634, 32'd4183, 32'd7919},
{32'd2570, 32'd3641, 32'd15166, -32'd1687},
{32'd772, -32'd4764, -32'd4670, -32'd2922},
{32'd793, -32'd16107, 32'd8820, 32'd4560},
{32'd1625, 32'd9924, 32'd2240, -32'd8926},
{32'd3046, -32'd4441, 32'd1393, 32'd6144},
{32'd4228, -32'd16654, 32'd7446, 32'd4628},
{32'd3818, 32'd14308, 32'd13098, -32'd5662},
{32'd4940, -32'd6852, -32'd9357, -32'd1086},
{-32'd223, 32'd8057, 32'd4430, 32'd7250},
{-32'd7727, -32'd11184, 32'd1689, 32'd7841},
{-32'd7771, 32'd1095, 32'd3741, -32'd5990},
{32'd11291, -32'd3373, 32'd7096, 32'd6867},
{-32'd7225, -32'd14453, 32'd12194, 32'd4870},
{32'd5945, -32'd10467, -32'd2738, 32'd7107},
{-32'd8800, 32'd2215, -32'd3375, 32'd6326},
{32'd3459, -32'd127, -32'd5736, 32'd13998},
{32'd9050, -32'd10919, 32'd1403, 32'd1192},
{-32'd3455, 32'd8619, 32'd7608, -32'd2200},
{32'd9532, -32'd1332, -32'd10980, -32'd6371},
{-32'd4653, -32'd12956, -32'd938, -32'd18714},
{32'd10190, 32'd1263, -32'd5801, -32'd577},
{32'd2256, 32'd305, 32'd4762, 32'd122},
{-32'd2885, -32'd11962, 32'd728, 32'd16545},
{-32'd4246, 32'd9875, -32'd8995, 32'd4111},
{-32'd3689, 32'd5086, -32'd1321, -32'd10622},
{-32'd643, 32'd8087, -32'd8913, 32'd535},
{32'd448, -32'd21985, 32'd10184, -32'd10176},
{32'd3983, 32'd1869, 32'd734, -32'd2282},
{32'd20867, -32'd3962, 32'd6, 32'd5327},
{-32'd1503, -32'd8312, 32'd2393, -32'd2707},
{32'd3897, 32'd1322, 32'd8217, 32'd5993},
{32'd1782, 32'd1994, 32'd3666, -32'd2815},
{32'd7776, -32'd12563, 32'd18403, 32'd10818},
{-32'd1622, 32'd1581, -32'd4974, 32'd6330},
{-32'd5066, 32'd8672, 32'd2473, -32'd2995},
{-32'd4823, 32'd65, -32'd6194, -32'd2560},
{32'd4314, -32'd7823, -32'd774, 32'd2264},
{32'd4358, 32'd16116, 32'd5049, 32'd10179},
{-32'd1033, 32'd8232, -32'd6053, 32'd1288},
{32'd554, -32'd1417, -32'd2292, 32'd7025},
{-32'd301, 32'd8814, -32'd1736, -32'd1474},
{32'd3285, -32'd9471, -32'd4636, 32'd10303},
{-32'd5634, 32'd6818, 32'd6015, -32'd1070},
{32'd10014, 32'd1321, 32'd5329, 32'd16573},
{-32'd1294, 32'd4112, -32'd8634, 32'd4960},
{32'd8238, 32'd16124, 32'd6354, -32'd578},
{32'd452, -32'd14771, 32'd696, -32'd5582},
{32'd1856, -32'd4418, -32'd6842, 32'd3041},
{32'd8750, -32'd3796, -32'd2362, -32'd3428},
{32'd5366, 32'd8101, -32'd2271, -32'd683},
{-32'd5131, 32'd12861, -32'd3025, 32'd3924},
{-32'd3740, -32'd33, -32'd5404, 32'd10334},
{32'd1312, -32'd22295, 32'd5426, -32'd3200},
{32'd698, 32'd1668, -32'd11679, 32'd5777},
{32'd6863, -32'd9601, -32'd4284, -32'd9337},
{32'd6875, 32'd15736, 32'd1172, 32'd324},
{32'd3921, 32'd19021, -32'd13390, 32'd1593},
{-32'd6586, -32'd5825, -32'd10458, -32'd270},
{32'd2807, -32'd2093, 32'd5645, -32'd6554},
{-32'd813, -32'd1754, -32'd3406, -32'd8121},
{32'd3887, 32'd15711, 32'd290, -32'd1881},
{-32'd6539, 32'd8740, -32'd11744, -32'd169},
{-32'd476, 32'd10685, -32'd4919, 32'd7515},
{32'd724, 32'd2817, 32'd10944, -32'd2102},
{-32'd2550, 32'd9618, 32'd1019, 32'd11290},
{32'd5648, -32'd20775, 32'd1756, -32'd1446},
{-32'd5716, 32'd1454, -32'd6519, 32'd5943},
{32'd2573, 32'd8077, 32'd2651, 32'd451},
{32'd664, 32'd16442, -32'd3311, -32'd1294},
{-32'd2691, 32'd3739, 32'd6837, -32'd6092},
{-32'd8965, 32'd3893, 32'd2819, -32'd773},
{32'd2728, -32'd66, -32'd1780, -32'd3649},
{32'd968, 32'd10289, 32'd4322, -32'd2696},
{32'd6983, 32'd9763, 32'd2243, -32'd3428},
{-32'd4633, -32'd3064, 32'd2303, -32'd3604},
{-32'd6476, -32'd1543, 32'd7255, -32'd12560},
{32'd13340, 32'd3078, -32'd1123, -32'd1282},
{32'd8037, -32'd2538, 32'd1384, 32'd6285},
{32'd537, 32'd3000, 32'd491, 32'd6883},
{-32'd3716, -32'd6794, -32'd4865, 32'd240},
{32'd3417, 32'd14742, -32'd5862, -32'd5952},
{32'd3796, -32'd8468, 32'd1625, 32'd1477},
{-32'd12893, -32'd1210, -32'd9213, 32'd2363},
{-32'd6289, -32'd6545, -32'd4772, 32'd1462},
{-32'd3256, -32'd12686, -32'd5135, -32'd15870},
{32'd9274, 32'd314, -32'd6527, 32'd5506},
{-32'd10184, -32'd4886, -32'd13884, -32'd5382},
{-32'd163, -32'd6979, 32'd6018, 32'd7998},
{-32'd8923, -32'd13273, 32'd14899, -32'd10700},
{-32'd2007, -32'd4391, 32'd3835, 32'd7908},
{-32'd5254, -32'd4737, -32'd1665, -32'd450},
{-32'd6616, -32'd7822, 32'd14185, 32'd3613},
{32'd1377, -32'd11593, 32'd504, -32'd5607},
{-32'd1041, -32'd6161, 32'd5626, -32'd6425},
{32'd4304, -32'd7361, 32'd11990, -32'd2610},
{32'd3441, 32'd12429, -32'd484, 32'd6407},
{32'd5953, -32'd15009, -32'd98, 32'd3824},
{-32'd144, 32'd18892, -32'd6744, 32'd3461},
{32'd3365, 32'd17674, 32'd3859, 32'd7689},
{-32'd70, -32'd5603, -32'd213, -32'd1130},
{32'd5196, 32'd6490, -32'd4076, -32'd5618},
{-32'd1401, -32'd4732, 32'd12054, 32'd10545},
{32'd234, -32'd6079, 32'd2280, -32'd5170},
{-32'd4280, -32'd15780, 32'd10248, 32'd3816},
{32'd1970, -32'd20187, 32'd6188, 32'd9740},
{-32'd11921, 32'd10932, 32'd3212, -32'd6771},
{-32'd3304, -32'd2512, 32'd6569, -32'd483},
{32'd1375, -32'd12749, 32'd8377, 32'd1043},
{-32'd2079, -32'd3285, 32'd6773, -32'd3892},
{-32'd6448, 32'd8118, -32'd8680, 32'd10160},
{32'd6828, 32'd22173, -32'd217, 32'd18465},
{32'd1885, 32'd8061, -32'd4694, 32'd9748},
{32'd1162, 32'd1231, -32'd3695, 32'd5483},
{32'd1952, -32'd9187, 32'd5957, -32'd5897},
{-32'd383, 32'd11192, -32'd718, 32'd5245},
{32'd844, 32'd3471, -32'd9985, 32'd624},
{32'd2643, -32'd4887, -32'd5500, -32'd9472},
{-32'd9040, 32'd17107, 32'd7835, -32'd6966},
{-32'd3448, 32'd4828, 32'd833, -32'd2933},
{-32'd1586, -32'd17612, -32'd9951, -32'd2189},
{-32'd1285, 32'd3379, 32'd3362, 32'd5626},
{32'd9215, -32'd16562, 32'd11017, -32'd1571},
{-32'd804, -32'd575, 32'd1905, -32'd9779},
{-32'd3450, -32'd18803, 32'd4797, 32'd5330},
{32'd10436, 32'd2593, 32'd1782, 32'd13713},
{32'd5415, -32'd19834, 32'd7919, -32'd5864},
{-32'd4430, 32'd1046, 32'd9625, -32'd2802},
{-32'd427, -32'd10106, -32'd14759, -32'd1945},
{-32'd856, -32'd1223, -32'd750, 32'd5671},
{-32'd6844, 32'd12885, -32'd9391, 32'd945},
{32'd898, 32'd6269, 32'd616, 32'd7414},
{-32'd2479, 32'd11871, 32'd4731, 32'd8166},
{32'd756, -32'd6560, -32'd1990, -32'd5678},
{32'd3847, -32'd1617, 32'd4364, -32'd6067},
{-32'd1236, 32'd188, -32'd4749, 32'd2320},
{32'd10086, 32'd5875, 32'd3363, 32'd6810},
{32'd7229, 32'd15332, 32'd3195, -32'd5413},
{-32'd10740, 32'd7652, -32'd3803, -32'd9409},
{-32'd4309, 32'd19756, -32'd2355, -32'd2444},
{-32'd91, -32'd6430, 32'd439, -32'd6112},
{32'd11212, 32'd23307, -32'd6796, 32'd1886},
{32'd2420, 32'd21135, 32'd5540, -32'd4125},
{32'd4222, 32'd8530, -32'd2988, -32'd3824},
{32'd3972, -32'd4254, 32'd3405, 32'd7953},
{-32'd5250, -32'd4850, -32'd3728, 32'd6137},
{32'd3425, 32'd3883, 32'd4287, -32'd11866},
{32'd1284, 32'd14820, 32'd9410, -32'd6560},
{32'd9913, -32'd2696, 32'd3780, -32'd2454},
{32'd6030, -32'd4103, 32'd17809, -32'd11467},
{32'd6052, 32'd8893, 32'd2161, 32'd4887},
{-32'd4427, -32'd1071, -32'd934, -32'd10594},
{-32'd3322, 32'd6204, 32'd7953, 32'd13540},
{-32'd667, -32'd244, -32'd7136, -32'd6611},
{32'd449, 32'd1543, -32'd2416, -32'd5320},
{-32'd5484, -32'd13177, -32'd2678, 32'd3270},
{-32'd5846, 32'd4678, -32'd3219, 32'd6583},
{-32'd5227, -32'd542, -32'd4135, -32'd2462},
{-32'd10261, -32'd1141, 32'd3792, 32'd2816},
{32'd525, 32'd11418, 32'd5443, 32'd3297},
{32'd1057, -32'd24677, 32'd9965, 32'd7868},
{-32'd2282, -32'd12768, -32'd2278, -32'd12162},
{32'd2506, -32'd6535, 32'd4194, -32'd3774},
{32'd124, 32'd7102, -32'd1739, -32'd11},
{-32'd2500, -32'd21779, -32'd3356, 32'd13178},
{-32'd2146, 32'd4922, 32'd4779, -32'd14435},
{32'd1347, -32'd12124, -32'd4456, -32'd4366},
{32'd7663, -32'd12374, 32'd9710, 32'd3544},
{32'd349, 32'd4694, -32'd608, 32'd2326},
{32'd5648, 32'd1119, 32'd3687, 32'd7785},
{-32'd2972, 32'd17593, 32'd2940, 32'd8535},
{-32'd7092, 32'd4479, -32'd2405, -32'd1573},
{-32'd7128, -32'd6716, -32'd1445, 32'd1292},
{32'd5360, -32'd2727, -32'd3226, 32'd10756},
{32'd1562, 32'd8195, -32'd3061, -32'd1313},
{-32'd1743, 32'd10612, -32'd2200, -32'd1854},
{32'd6878, -32'd6430, -32'd7467, 32'd4382},
{-32'd10469, 32'd1393, 32'd1611, 32'd335},
{32'd754, -32'd8939, -32'd11708, -32'd6043},
{32'd1227, -32'd6009, -32'd10040, 32'd7072},
{-32'd1647, -32'd882, -32'd12873, -32'd3572},
{-32'd1399, -32'd22818, 32'd9132, 32'd9488},
{32'd11364, -32'd9534, -32'd4798, -32'd1262},
{32'd5108, 32'd1652, 32'd1427, 32'd2756},
{-32'd221, 32'd9311, -32'd1731, -32'd2474},
{-32'd5042, 32'd14579, 32'd2131, 32'd701},
{-32'd4892, 32'd1333, 32'd6692, -32'd11198},
{-32'd11234, -32'd4171, -32'd16201, -32'd4350},
{-32'd8273, 32'd10350, 32'd2506, 32'd4769},
{32'd6083, -32'd9051, 32'd8825, -32'd4432},
{32'd5365, -32'd3488, 32'd13062, 32'd3773},
{-32'd711, -32'd9637, -32'd4603, 32'd4924},
{-32'd3117, -32'd15531, -32'd5578, -32'd9817}
},
{{-32'd175, -32'd9906, -32'd3455, 32'd2205},
{32'd1153, 32'd9120, -32'd10060, 32'd4880},
{-32'd9105, -32'd11063, -32'd3859, -32'd12322},
{-32'd5013, 32'd7593, 32'd8578, 32'd1993},
{32'd10956, -32'd9697, 32'd14287, 32'd6341},
{-32'd8111, 32'd192, 32'd2901, -32'd7570},
{-32'd9649, 32'd14409, 32'd10965, 32'd13072},
{-32'd9086, 32'd4252, -32'd13442, -32'd4649},
{-32'd18217, -32'd3, 32'd1191, 32'd4574},
{-32'd3952, 32'd2966, 32'd5048, 32'd10971},
{32'd5821, -32'd7005, -32'd5120, 32'd9522},
{-32'd7179, -32'd7102, -32'd5249, -32'd6050},
{32'd883, 32'd19009, -32'd11881, -32'd8190},
{32'd337, -32'd7497, -32'd254, 32'd6607},
{32'd1045, 32'd2402, 32'd1981, -32'd10475},
{32'd10191, -32'd7235, -32'd6708, -32'd2171},
{32'd345, -32'd533, 32'd2191, 32'd1463},
{-32'd1507, -32'd5237, -32'd3750, 32'd9629},
{-32'd8470, -32'd11666, -32'd7930, -32'd3508},
{-32'd16, -32'd5992, -32'd15561, 32'd14564},
{-32'd7763, 32'd7266, 32'd5054, 32'd3184},
{32'd1485, -32'd3930, 32'd201, 32'd3480},
{-32'd3237, 32'd6818, -32'd13239, -32'd9007},
{32'd7106, -32'd1423, -32'd4622, 32'd3655},
{-32'd1245, 32'd668, -32'd7926, -32'd2983},
{-32'd5393, -32'd11103, 32'd8975, -32'd7273},
{-32'd11280, 32'd1813, -32'd12459, 32'd1026},
{32'd905, -32'd3061, 32'd4348, 32'd6060},
{32'd986, 32'd4816, 32'd7045, 32'd6779},
{32'd6045, 32'd7342, 32'd2176, 32'd9430},
{32'd22487, 32'd2092, -32'd7607, -32'd3586},
{-32'd3897, 32'd1673, -32'd3688, -32'd3076},
{-32'd2973, 32'd580, -32'd1455, -32'd3001},
{32'd11493, -32'd14763, -32'd750, -32'd1982},
{-32'd2538, 32'd8604, 32'd3606, 32'd9561},
{-32'd8025, 32'd3906, -32'd4220, 32'd2763},
{32'd4737, -32'd1231, 32'd12154, 32'd7043},
{-32'd17654, -32'd9021, 32'd25091, 32'd10864},
{32'd3590, 32'd2987, -32'd9872, -32'd13177},
{-32'd13553, 32'd6394, -32'd3285, -32'd642},
{-32'd3063, -32'd4073, 32'd4680, 32'd2581},
{32'd4712, 32'd6651, -32'd11594, 32'd17457},
{32'd4122, -32'd7658, 32'd1033, 32'd14508},
{32'd15583, 32'd8744, -32'd10506, -32'd13408},
{32'd4451, -32'd6547, -32'd14588, -32'd8886},
{32'd10521, -32'd6447, 32'd725, 32'd8660},
{-32'd7081, 32'd6826, -32'd3977, 32'd18986},
{32'd587, -32'd4099, -32'd3452, -32'd2643},
{-32'd5084, 32'd2312, 32'd1411, 32'd372},
{-32'd11349, 32'd4869, 32'd5973, -32'd688},
{32'd4695, 32'd5322, -32'd6609, 32'd5684},
{-32'd8204, 32'd10810, -32'd8576, -32'd14220},
{32'd5847, -32'd9724, -32'd6464, 32'd3776},
{32'd9791, -32'd5831, 32'd573, -32'd272},
{32'd16960, 32'd6782, -32'd5269, 32'd1035},
{32'd8169, 32'd8075, -32'd1427, -32'd8196},
{32'd2171, 32'd5248, 32'd12397, -32'd4684},
{32'd17996, -32'd5880, -32'd4172, -32'd152},
{32'd11962, -32'd8775, -32'd6523, -32'd3791},
{-32'd18440, 32'd9886, -32'd2623, -32'd6230},
{32'd2206, 32'd15089, 32'd7026, 32'd6441},
{-32'd7182, 32'd5213, 32'd8065, -32'd6639},
{32'd5013, -32'd7398, -32'd6130, 32'd1853},
{-32'd1866, 32'd9986, 32'd1296, -32'd4369},
{32'd9595, -32'd7865, 32'd2071, -32'd8638},
{-32'd6388, 32'd11606, -32'd6585, 32'd12939},
{-32'd515, -32'd1099, 32'd7995, -32'd4863},
{32'd3123, 32'd6768, -32'd16386, 32'd1057},
{32'd82, -32'd5530, -32'd17638, -32'd7645},
{-32'd6452, -32'd5355, -32'd1428, -32'd1914},
{32'd7443, 32'd3592, -32'd1623, -32'd9882},
{32'd8375, 32'd14293, 32'd448, 32'd11620},
{32'd4960, -32'd2625, -32'd12171, 32'd695},
{-32'd6515, 32'd6582, -32'd2654, 32'd6035},
{-32'd5191, 32'd1674, 32'd9664, 32'd7496},
{32'd6901, 32'd1597, 32'd790, -32'd9297},
{-32'd231, -32'd3907, 32'd9602, -32'd3457},
{-32'd433, -32'd3376, 32'd918, -32'd6929},
{32'd4194, 32'd12435, -32'd889, 32'd13302},
{32'd4495, -32'd8171, 32'd12369, 32'd1522},
{-32'd4451, -32'd3934, -32'd9114, -32'd1847},
{32'd2080, -32'd6371, -32'd5603, 32'd8439},
{-32'd3154, 32'd4917, 32'd47, -32'd5045},
{32'd5390, -32'd2231, 32'd5733, -32'd117},
{32'd4949, -32'd7741, 32'd864, -32'd2627},
{32'd17537, 32'd7644, -32'd7040, -32'd5862},
{32'd1829, -32'd8479, -32'd2589, 32'd4440},
{32'd5994, -32'd3860, -32'd9525, -32'd3969},
{32'd16666, -32'd9446, 32'd4353, -32'd6608},
{32'd1812, -32'd128, 32'd3007, -32'd9942},
{-32'd4904, 32'd4329, -32'd6555, 32'd8379},
{-32'd6564, 32'd8962, -32'd4569, 32'd4142},
{-32'd501, -32'd22485, -32'd1022, 32'd4146},
{32'd5848, 32'd7503, -32'd6449, 32'd8714},
{-32'd1092, 32'd3320, 32'd5367, 32'd7437},
{-32'd784, -32'd8499, 32'd4054, 32'd981},
{-32'd3757, -32'd1462, 32'd434, 32'd5730},
{-32'd10401, 32'd1873, 32'd442, -32'd9365},
{32'd4011, 32'd4512, 32'd809, -32'd2811},
{-32'd11741, -32'd2932, 32'd9966, 32'd684},
{-32'd3957, -32'd4510, 32'd188, -32'd10281},
{32'd2206, -32'd4367, -32'd20614, 32'd3430},
{32'd4697, 32'd1565, 32'd19326, 32'd3162},
{-32'd2906, -32'd415, 32'd10283, -32'd1132},
{32'd384, -32'd483, -32'd2783, 32'd3965},
{32'd5962, -32'd509, -32'd4626, 32'd9048},
{-32'd8456, -32'd6977, 32'd3435, 32'd8350},
{-32'd12680, 32'd1391, -32'd6531, -32'd4192},
{32'd7972, 32'd4475, -32'd9597, 32'd2323},
{32'd4777, -32'd216, -32'd4080, -32'd6279},
{32'd12980, -32'd14868, 32'd438, -32'd1907},
{32'd5101, -32'd11666, 32'd5392, 32'd6800},
{32'd1592, 32'd12886, 32'd2358, 32'd15042},
{32'd10415, 32'd1873, 32'd3970, 32'd4767},
{32'd1085, -32'd13743, -32'd4369, 32'd3090},
{-32'd3634, 32'd7589, -32'd7413, 32'd13903},
{-32'd5089, -32'd1392, -32'd6536, -32'd10041},
{-32'd13492, 32'd17265, 32'd4241, 32'd3343},
{32'd6116, -32'd1354, 32'd6977, 32'd9696},
{-32'd2594, 32'd5572, 32'd7316, 32'd6591},
{-32'd5783, 32'd8365, -32'd18035, -32'd1039},
{-32'd3723, -32'd11648, 32'd5595, -32'd5812},
{-32'd2831, -32'd4022, -32'd3311, -32'd2950},
{-32'd6353, -32'd7605, 32'd13979, 32'd9569},
{32'd3878, -32'd12946, 32'd2385, -32'd168},
{-32'd3859, 32'd10538, 32'd454, 32'd1184},
{-32'd1197, -32'd1676, 32'd1835, -32'd14212},
{32'd13642, -32'd12953, -32'd7504, -32'd7111},
{32'd3074, -32'd6279, 32'd4506, -32'd1851},
{-32'd9833, -32'd5960, -32'd3641, -32'd3013},
{-32'd5457, 32'd3100, -32'd3690, 32'd1057},
{-32'd6765, -32'd4008, -32'd10467, 32'd4770},
{32'd12833, -32'd14706, -32'd1857, -32'd717},
{-32'd11964, 32'd11410, 32'd2464, -32'd7104},
{32'd3132, 32'd3854, -32'd14341, 32'd5733},
{32'd12583, 32'd6008, 32'd5626, 32'd9483},
{32'd10159, 32'd4765, -32'd7139, 32'd21930},
{-32'd574, -32'd19525, 32'd176, -32'd29},
{32'd3786, 32'd9104, 32'd10913, 32'd4027},
{-32'd1281, -32'd1041, -32'd445, 32'd2878},
{-32'd6369, -32'd7195, 32'd2838, 32'd2097},
{32'd4169, 32'd715, -32'd4983, 32'd3128},
{-32'd1481, -32'd2785, -32'd845, -32'd3170},
{32'd13075, -32'd493, -32'd9800, -32'd3972},
{32'd2156, 32'd1754, 32'd2454, -32'd1521},
{-32'd5067, 32'd3149, 32'd10670, -32'd455},
{-32'd2575, -32'd15486, -32'd476, -32'd1470},
{32'd3334, -32'd8345, 32'd7792, -32'd7888},
{-32'd8312, 32'd20148, -32'd1488, -32'd597},
{-32'd197, -32'd9404, -32'd8435, -32'd8520},
{32'd6732, -32'd14544, 32'd4080, -32'd6279},
{32'd3369, -32'd5380, 32'd8432, 32'd10754},
{32'd1591, -32'd12240, 32'd2832, 32'd4230},
{32'd5950, 32'd5461, -32'd7585, -32'd804},
{32'd8010, -32'd2873, -32'd2024, 32'd4764},
{32'd14269, -32'd6704, 32'd8245, -32'd3312},
{-32'd5322, -32'd8279, -32'd16947, 32'd12373},
{32'd6859, -32'd1445, 32'd12400, -32'd2869},
{-32'd7884, -32'd847, 32'd3849, 32'd8509},
{-32'd3541, 32'd3793, -32'd2997, 32'd8073},
{-32'd2175, 32'd1729, -32'd743, 32'd6784},
{32'd3731, 32'd1761, -32'd7488, -32'd15108},
{-32'd912, -32'd17673, 32'd3607, 32'd7187},
{-32'd1863, -32'd1321, 32'd8151, -32'd3252},
{-32'd12957, 32'd15684, 32'd8510, -32'd4920},
{-32'd7309, 32'd14216, -32'd5131, 32'd3294},
{-32'd3753, 32'd7709, -32'd2415, -32'd494},
{32'd18094, -32'd6905, -32'd4171, 32'd859},
{32'd13807, 32'd4349, 32'd7191, 32'd3079},
{-32'd6563, -32'd5019, -32'd1200, -32'd21939},
{-32'd13237, 32'd7799, 32'd7480, -32'd4754},
{-32'd20879, 32'd2455, 32'd8413, 32'd9565},
{-32'd83, 32'd10861, 32'd633, 32'd8011},
{-32'd21907, -32'd4455, 32'd796, 32'd1174},
{-32'd2896, 32'd10851, 32'd3696, -32'd1758},
{32'd14624, -32'd6594, -32'd6517, -32'd9359},
{-32'd1237, -32'd2879, 32'd15065, -32'd8905},
{-32'd14706, 32'd10750, 32'd7647, 32'd1372},
{-32'd9524, -32'd5604, 32'd2197, 32'd9970},
{32'd6942, 32'd68, -32'd2063, -32'd9153},
{-32'd1196, -32'd3561, -32'd2337, 32'd985},
{32'd12748, -32'd13009, -32'd9956, -32'd4203},
{32'd1953, 32'd6611, -32'd11370, -32'd9303},
{32'd2997, 32'd5286, 32'd6898, 32'd518},
{-32'd4681, -32'd16714, -32'd5200, 32'd7212},
{32'd458, 32'd8722, 32'd4449, 32'd386},
{-32'd10558, 32'd6251, -32'd1566, 32'd6949},
{-32'd5134, -32'd3595, 32'd7183, 32'd6615},
{32'd6942, 32'd4308, 32'd9627, 32'd13479},
{32'd12559, -32'd6843, 32'd2387, 32'd2601},
{32'd14485, 32'd13056, -32'd870, 32'd5851},
{32'd1783, -32'd3626, -32'd19976, -32'd3614},
{-32'd2667, 32'd8639, -32'd3063, -32'd11434},
{32'd359, 32'd6023, -32'd4134, 32'd5917},
{-32'd14816, 32'd7127, 32'd2677, -32'd3632},
{32'd2816, -32'd17754, -32'd1075, -32'd10964},
{-32'd8105, -32'd2871, 32'd14210, -32'd3494},
{32'd346, -32'd2446, -32'd120, -32'd6012},
{32'd414, -32'd14918, -32'd13212, -32'd2017},
{-32'd2298, -32'd6930, 32'd3386, 32'd2606},
{32'd6029, -32'd7521, -32'd1800, -32'd6622},
{-32'd1808, 32'd3585, -32'd10235, -32'd4987},
{32'd12440, -32'd8064, -32'd2731, 32'd9140},
{-32'd7633, -32'd5192, 32'd15470, 32'd20563},
{-32'd4790, 32'd271, -32'd6865, 32'd1712},
{32'd6057, -32'd10463, 32'd3837, 32'd4457},
{-32'd4901, 32'd1181, 32'd5399, 32'd2210},
{32'd4321, 32'd2851, 32'd1522, -32'd10708},
{32'd15364, -32'd6802, -32'd12171, -32'd5679},
{32'd4041, -32'd8823, 32'd157, -32'd5207},
{32'd14072, 32'd1283, 32'd406, -32'd9550},
{-32'd4831, 32'd3777, 32'd264, 32'd3516},
{32'd1018, -32'd7097, -32'd6575, -32'd7187},
{-32'd17620, -32'd1259, 32'd2968, -32'd2253},
{32'd4597, -32'd9635, -32'd6959, 32'd4036},
{-32'd1229, 32'd8890, -32'd12681, -32'd7696},
{-32'd6764, 32'd14527, -32'd6160, 32'd10394},
{-32'd2747, 32'd1992, 32'd9815, -32'd5543},
{-32'd16526, 32'd1418, 32'd7031, 32'd2633},
{-32'd8048, -32'd333, 32'd4159, -32'd4832},
{32'd11065, -32'd4592, -32'd10024, 32'd4109},
{-32'd9082, 32'd5231, 32'd3396, 32'd14621},
{32'd10534, 32'd5083, 32'd11780, 32'd4421},
{32'd4344, -32'd167, 32'd2297, -32'd3169},
{32'd7568, -32'd1090, -32'd7236, -32'd12572},
{32'd439, 32'd6837, -32'd606, 32'd8561},
{-32'd2414, -32'd607, 32'd2919, 32'd8456},
{-32'd4793, 32'd1116, -32'd11497, 32'd2359},
{-32'd8653, -32'd7167, -32'd3656, 32'd2129},
{32'd19075, 32'd10776, 32'd650, -32'd2356},
{-32'd5720, -32'd13291, -32'd6141, -32'd3931},
{32'd2584, -32'd14445, 32'd1023, -32'd6579},
{-32'd11555, 32'd1039, -32'd337, -32'd1956},
{32'd16423, 32'd1278, -32'd9876, 32'd1525},
{32'd2792, 32'd3155, -32'd9944, -32'd1317},
{32'd7005, 32'd5753, 32'd17423, 32'd5222},
{-32'd8035, -32'd2571, -32'd6278, 32'd4686},
{-32'd3974, 32'd11693, -32'd1745, 32'd8701},
{-32'd975, 32'd1538, 32'd2125, -32'd2007},
{32'd4765, 32'd5410, -32'd9728, -32'd8040},
{-32'd3475, -32'd2935, 32'd4396, 32'd6541},
{32'd7252, -32'd6999, 32'd956, 32'd7899},
{32'd7358, -32'd7895, -32'd3967, -32'd10103},
{-32'd903, -32'd2879, 32'd11838, 32'd2598},
{32'd3780, 32'd8961, 32'd8204, 32'd4146},
{-32'd2682, -32'd4416, -32'd1891, -32'd11045},
{32'd1441, 32'd5384, 32'd3760, 32'd5267},
{-32'd18406, 32'd6152, 32'd5882, 32'd2051},
{32'd1088, -32'd3189, 32'd1048, -32'd3797},
{-32'd9355, 32'd6187, 32'd2704, -32'd5777},
{32'd17633, 32'd7774, -32'd1846, -32'd200},
{32'd457, -32'd6776, 32'd1178, -32'd7788},
{32'd2936, -32'd4746, 32'd4820, 32'd11250},
{32'd3425, 32'd7748, -32'd13843, 32'd1291},
{32'd9414, -32'd3611, 32'd114, 32'd5131},
{-32'd745, 32'd346, 32'd4869, 32'd12484},
{32'd9821, 32'd6545, -32'd4090, -32'd11661},
{-32'd1577, -32'd3530, 32'd7839, -32'd4984},
{32'd2918, -32'd15867, 32'd4278, -32'd5312},
{-32'd7287, -32'd5259, 32'd6424, 32'd4140},
{-32'd13534, 32'd20149, 32'd6224, 32'd230},
{32'd11724, 32'd1185, 32'd5280, -32'd12591},
{-32'd10036, -32'd117, -32'd1191, 32'd3311},
{-32'd3199, 32'd6786, -32'd4190, -32'd1199},
{-32'd2406, 32'd5519, 32'd1135, -32'd4408},
{32'd2877, 32'd8179, -32'd7758, -32'd158},
{32'd3282, -32'd9378, 32'd10544, -32'd14311},
{32'd11549, -32'd7322, -32'd2607, -32'd2870},
{32'd12203, 32'd2620, -32'd7258, -32'd507},
{32'd3216, 32'd13997, 32'd10258, -32'd7670},
{32'd1514, 32'd11451, 32'd7903, 32'd2600},
{-32'd5828, 32'd6142, 32'd4843, -32'd6726},
{32'd20239, -32'd981, 32'd5059, -32'd7278},
{-32'd5790, 32'd8592, -32'd7576, 32'd1628},
{32'd3629, -32'd2870, -32'd14934, -32'd11324},
{-32'd5527, 32'd8185, -32'd985, 32'd887},
{-32'd2196, 32'd8265, 32'd1745, 32'd10573},
{-32'd14330, -32'd1956, -32'd861, -32'd11005},
{32'd8751, -32'd11912, -32'd5177, -32'd14465},
{32'd1921, 32'd4366, 32'd1498, 32'd3141},
{-32'd12040, -32'd2689, 32'd373, 32'd4822},
{-32'd3906, -32'd2686, 32'd6505, 32'd16572},
{32'd7858, -32'd2837, 32'd7703, -32'd4499},
{-32'd12214, 32'd9319, -32'd3584, -32'd1233},
{-32'd13532, 32'd6113, -32'd12106, -32'd2360},
{32'd1325, -32'd8024, -32'd9744, -32'd4579},
{-32'd770, -32'd9359, 32'd2696, 32'd13711},
{32'd7666, -32'd4866, -32'd165, -32'd1600},
{-32'd6579, 32'd8769, 32'd3552, 32'd14159},
{32'd10085, -32'd7366, -32'd7027, 32'd3325},
{32'd3789, -32'd3093, -32'd4853, -32'd14078},
{-32'd1136, -32'd886, -32'd1, 32'd8196},
{-32'd3976, -32'd5057, 32'd1573, -32'd7578},
{-32'd9879, -32'd1189, -32'd4642, 32'd4861},
{-32'd2771, 32'd1839, -32'd5377, -32'd16543},
{32'd6873, -32'd3933, 32'd1029, -32'd6680},
{32'd9123, 32'd3263, -32'd3789, -32'd3231},
{32'd6164, -32'd8605, -32'd5628, 32'd3021},
{-32'd4961, 32'd9446, -32'd10879, 32'd1363},
{32'd1506, -32'd5517, 32'd1916, 32'd3334}
},
{{32'd10369, 32'd10072, 32'd7188, -32'd1199},
{-32'd776, -32'd6733, -32'd469, -32'd5446},
{32'd17957, -32'd382, -32'd3026, 32'd2623},
{32'd9978, 32'd5304, 32'd6967, 32'd2162},
{32'd3595, -32'd2236, 32'd10604, 32'd1693},
{32'd7179, -32'd10170, 32'd6227, -32'd5082},
{-32'd3963, 32'd4565, -32'd227, -32'd2541},
{-32'd5554, 32'd1927, -32'd3494, 32'd648},
{32'd5673, 32'd7028, 32'd8743, -32'd5563},
{32'd9285, 32'd15822, 32'd9816, 32'd5229},
{32'd16530, -32'd6706, 32'd4209, -32'd99},
{-32'd2520, 32'd566, -32'd3920, -32'd5209},
{32'd3503, 32'd7631, 32'd8346, -32'd7514},
{-32'd2480, 32'd1663, -32'd9847, -32'd9315},
{-32'd179, -32'd6247, 32'd478, 32'd6089},
{32'd2385, -32'd404, 32'd5312, -32'd1476},
{32'd9095, 32'd11686, 32'd16226, 32'd497},
{-32'd1849, 32'd11678, -32'd3476, 32'd7212},
{-32'd363, 32'd475, -32'd11198, -32'd4446},
{32'd6627, 32'd932, 32'd12372, -32'd4814},
{-32'd1707, 32'd6768, 32'd7173, 32'd2793},
{32'd4839, -32'd3185, -32'd1972, -32'd8992},
{32'd315, 32'd1976, 32'd4553, -32'd7477},
{32'd436, -32'd10226, -32'd12088, -32'd10689},
{32'd2346, -32'd2152, 32'd18254, 32'd8245},
{-32'd4881, 32'd4077, -32'd7382, -32'd7295},
{32'd991, -32'd6622, 32'd5985, -32'd9438},
{-32'd1410, 32'd3029, -32'd12249, 32'd2416},
{32'd854, 32'd5192, 32'd15290, -32'd8464},
{-32'd14752, -32'd3671, -32'd3219, -32'd13691},
{32'd4096, -32'd4649, -32'd3067, 32'd593},
{-32'd9689, -32'd8056, -32'd10742, -32'd13220},
{32'd2614, 32'd7279, 32'd4755, 32'd1235},
{-32'd15739, 32'd3242, -32'd7985, 32'd1737},
{32'd2536, 32'd9846, 32'd9280, -32'd789},
{-32'd4291, -32'd6167, -32'd6687, -32'd655},
{32'd141, -32'd6626, -32'd1282, 32'd58},
{-32'd1443, 32'd4840, 32'd6486, 32'd2466},
{-32'd2578, 32'd10876, 32'd8314, -32'd353},
{32'd6306, 32'd2845, 32'd6902, 32'd4662},
{32'd8691, 32'd6009, 32'd9401, -32'd988},
{32'd775, 32'd4203, 32'd2770, -32'd5851},
{32'd11057, 32'd4288, 32'd1779, 32'd11014},
{-32'd1025, -32'd5143, -32'd4381, 32'd6015},
{-32'd3813, -32'd10217, -32'd6337, -32'd2950},
{-32'd5010, 32'd1536, 32'd126, 32'd1412},
{-32'd3192, -32'd9421, -32'd2939, 32'd2958},
{32'd922, 32'd1687, -32'd15652, -32'd5503},
{32'd11288, 32'd12029, 32'd17929, 32'd10267},
{32'd1876, -32'd5110, -32'd625, 32'd12496},
{-32'd7701, -32'd1296, 32'd6482, -32'd13590},
{-32'd6033, 32'd3627, -32'd4620, 32'd9383},
{-32'd1939, -32'd2819, -32'd7169, -32'd6109},
{32'd5192, -32'd3393, 32'd202, 32'd4687},
{32'd5856, 32'd14179, 32'd6015, 32'd1930},
{32'd4978, -32'd2260, 32'd1194, -32'd10487},
{32'd6751, 32'd16561, 32'd6774, 32'd7509},
{-32'd17003, -32'd11095, -32'd10529, -32'd3659},
{-32'd5324, -32'd6812, -32'd7677, -32'd2915},
{-32'd17408, -32'd3105, -32'd6666, -32'd10621},
{-32'd16290, -32'd9679, -32'd11329, -32'd7590},
{32'd1225, 32'd7680, -32'd12384, 32'd7849},
{-32'd11570, -32'd6892, -32'd16667, -32'd10131},
{-32'd13358, -32'd3114, -32'd5379, 32'd10146},
{-32'd5057, 32'd6609, -32'd1465, 32'd7135},
{-32'd3591, 32'd1316, 32'd13949, 32'd2912},
{32'd507, -32'd700, 32'd7690, -32'd8511},
{-32'd10873, -32'd3431, -32'd7190, 32'd4389},
{-32'd1669, 32'd4032, 32'd1963, 32'd10742},
{-32'd7484, -32'd77, -32'd4699, -32'd2721},
{32'd13535, -32'd1123, 32'd868, 32'd10431},
{32'd2364, -32'd5844, -32'd6057, -32'd1865},
{-32'd8223, -32'd114, -32'd1061, 32'd7215},
{32'd7090, -32'd1957, 32'd21681, 32'd16605},
{-32'd116, 32'd7333, 32'd3195, -32'd2877},
{-32'd354, -32'd3714, 32'd4947, 32'd462},
{-32'd15, -32'd8153, -32'd10277, 32'd2969},
{-32'd11046, 32'd1643, -32'd1868, -32'd4576},
{-32'd814, 32'd2845, 32'd10699, 32'd6159},
{-32'd1161, 32'd4512, 32'd2980, 32'd3383},
{32'd5279, 32'd10243, 32'd8175, 32'd10758},
{32'd19395, 32'd2664, 32'd9540, 32'd17143},
{-32'd496, -32'd5790, -32'd2687, -32'd7920},
{32'd5795, 32'd9818, 32'd954, 32'd6952},
{-32'd18095, 32'd1565, 32'd1175, -32'd513},
{32'd2807, -32'd152, 32'd1513, 32'd120},
{-32'd200, 32'd3194, 32'd5300, -32'd7662},
{-32'd6457, -32'd6941, -32'd5524, 32'd4805},
{32'd5249, 32'd3899, 32'd11106, 32'd5856},
{32'd851, -32'd1893, -32'd16075, -32'd1617},
{32'd5270, -32'd2725, 32'd5089, 32'd7509},
{32'd2645, -32'd2276, -32'd568, -32'd4635},
{32'd2671, 32'd4930, 32'd10187, 32'd6558},
{-32'd10342, 32'd5586, 32'd8988, 32'd882},
{-32'd4535, 32'd5159, -32'd2346, 32'd7919},
{32'd9727, -32'd7851, -32'd2146, -32'd74},
{-32'd979, 32'd5755, 32'd1637, 32'd12898},
{-32'd8246, 32'd4917, -32'd2240, -32'd2069},
{32'd8616, -32'd6052, 32'd5909, -32'd4033},
{-32'd657, 32'd10705, -32'd351, 32'd3318},
{-32'd6300, 32'd10, 32'd6390, 32'd6166},
{32'd16394, -32'd1750, -32'd4600, 32'd4198},
{32'd3461, -32'd12954, -32'd6313, 32'd866},
{32'd14299, -32'd6098, 32'd8933, -32'd1161},
{32'd319, 32'd9380, 32'd12406, 32'd8059},
{-32'd2649, -32'd5213, -32'd2433, 32'd11335},
{-32'd4051, -32'd9456, -32'd2936, -32'd7993},
{32'd4055, -32'd3184, 32'd907, -32'd1992},
{32'd9675, 32'd321, 32'd7669, -32'd9020},
{32'd463, -32'd8100, -32'd10682, 32'd710},
{-32'd9378, 32'd676, -32'd5447, -32'd5546},
{-32'd4285, 32'd1089, -32'd7116, -32'd5820},
{32'd3934, 32'd8555, 32'd2870, 32'd5891},
{-32'd4966, -32'd7433, -32'd350, -32'd999},
{-32'd3649, -32'd3377, 32'd2223, -32'd9560},
{32'd2200, -32'd3044, 32'd1436, 32'd4217},
{-32'd5103, 32'd4133, 32'd4844, -32'd1644},
{-32'd5603, -32'd5263, 32'd518, 32'd462},
{-32'd2715, -32'd6398, -32'd3364, 32'd7876},
{-32'd4329, 32'd6202, 32'd6088, -32'd5030},
{32'd2782, 32'd3481, 32'd8135, 32'd14561},
{32'd1758, 32'd2617, -32'd11111, 32'd1732},
{-32'd4988, -32'd1300, -32'd1090, 32'd1561},
{32'd6872, -32'd10317, -32'd1499, -32'd2258},
{32'd6648, -32'd1941, -32'd585, 32'd7075},
{32'd4689, -32'd715, 32'd5407, -32'd7101},
{-32'd13261, -32'd3290, -32'd8340, 32'd201},
{32'd5933, 32'd6983, -32'd4756, 32'd12810},
{32'd3081, 32'd1115, -32'd10559, -32'd19679},
{32'd3843, 32'd728, -32'd1202, 32'd6681},
{-32'd2215, -32'd3823, 32'd11409, -32'd6643},
{-32'd14409, -32'd15984, 32'd3398, 32'd552},
{-32'd12520, -32'd7273, 32'd2117, 32'd5999},
{32'd11726, -32'd2205, 32'd6673, 32'd2872},
{32'd10447, -32'd5985, -32'd7499, -32'd4531},
{-32'd15386, 32'd5161, -32'd5439, 32'd7934},
{-32'd3195, 32'd2269, 32'd120, 32'd4112},
{32'd10127, -32'd8365, -32'd7795, -32'd3537},
{32'd1898, 32'd3143, 32'd845, 32'd2393},
{-32'd10039, 32'd3980, 32'd5110, 32'd4066},
{32'd2025, 32'd3644, -32'd8682, -32'd5374},
{-32'd9097, -32'd2542, -32'd7902, 32'd725},
{32'd2660, 32'd412, -32'd11385, 32'd3111},
{32'd9229, -32'd1373, 32'd3983, 32'd7},
{32'd1035, 32'd2986, -32'd9180, -32'd2113},
{32'd12888, 32'd7128, 32'd3388, 32'd5919},
{32'd6314, -32'd3785, -32'd1730, 32'd887},
{-32'd1162, -32'd6712, -32'd397, 32'd692},
{-32'd4816, 32'd2009, 32'd737, -32'd2436},
{32'd2992, -32'd15329, -32'd7106, 32'd1650},
{32'd2764, -32'd4616, -32'd9263, 32'd798},
{32'd7766, 32'd11, 32'd3791, 32'd1551},
{-32'd2417, -32'd2477, -32'd7685, -32'd3142},
{32'd9850, 32'd3298, 32'd4231, -32'd4861},
{32'd9803, -32'd10548, -32'd3663, 32'd3351},
{-32'd1010, 32'd3847, -32'd1466, -32'd4021},
{32'd13133, 32'd6530, 32'd2724, -32'd1901},
{32'd10987, 32'd465, 32'd11361, -32'd707},
{32'd5948, -32'd527, -32'd1090, -32'd11442},
{-32'd1979, 32'd4056, 32'd1450, 32'd887},
{32'd9866, -32'd10958, 32'd3249, -32'd14860},
{-32'd10130, 32'd5965, -32'd1110, -32'd3633},
{-32'd5702, -32'd7175, 32'd3143, -32'd11205},
{-32'd877, 32'd187, 32'd1641, 32'd10975},
{32'd11375, 32'd4648, 32'd12371, 32'd4933},
{-32'd10046, -32'd10466, 32'd3807, -32'd4223},
{-32'd16833, 32'd6696, 32'd6766, 32'd8985},
{-32'd1741, -32'd16828, -32'd2089, -32'd5322},
{-32'd6310, -32'd17094, -32'd5089, -32'd4393},
{-32'd5876, -32'd8012, -32'd8102, -32'd3928},
{32'd4341, 32'd2021, -32'd4924, 32'd2734},
{-32'd253, -32'd5950, -32'd5595, -32'd14156},
{32'd6797, 32'd9532, 32'd1109, -32'd1965},
{-32'd7185, -32'd1110, -32'd8558, -32'd5372},
{-32'd6713, 32'd13838, -32'd3089, -32'd2005},
{-32'd849, 32'd4502, -32'd1192, 32'd7473},
{-32'd881, 32'd10251, -32'd4652, 32'd12502},
{32'd6152, 32'd8916, 32'd3726, -32'd1106},
{32'd1648, 32'd4168, 32'd3992, 32'd11323},
{32'd1801, -32'd1940, -32'd3093, 32'd68},
{-32'd6452, -32'd11182, -32'd7332, 32'd3336},
{-32'd4964, -32'd3187, -32'd6802, 32'd8818},
{-32'd6084, -32'd1314, -32'd3126, -32'd6331},
{32'd3695, -32'd3844, -32'd3201, 32'd6742},
{-32'd7170, 32'd608, 32'd2894, 32'd7125},
{-32'd5103, 32'd6546, 32'd355, -32'd2456},
{-32'd2895, -32'd2524, -32'd3801, -32'd7054},
{32'd4223, -32'd318, -32'd3149, 32'd3259},
{-32'd10404, -32'd4214, 32'd6288, 32'd843},
{32'd2881, -32'd478, -32'd8592, -32'd4647},
{-32'd4619, 32'd338, 32'd10466, 32'd977},
{-32'd8584, -32'd11741, -32'd6144, -32'd441},
{32'd2864, -32'd5293, -32'd4014, -32'd1987},
{32'd2972, -32'd3462, 32'd3784, 32'd3661},
{32'd2591, -32'd909, -32'd1270, 32'd2594},
{32'd11024, 32'd1975, -32'd4486, -32'd9480},
{32'd2354, 32'd4866, -32'd14089, -32'd5112},
{32'd29774, 32'd5251, 32'd8572, -32'd1273},
{32'd6547, 32'd3236, -32'd1828, 32'd8035},
{32'd12038, -32'd967, 32'd8245, 32'd3954},
{32'd4487, -32'd8943, -32'd5544, -32'd1045},
{-32'd2908, -32'd4421, 32'd1152, -32'd8312},
{-32'd4500, 32'd3500, 32'd812, 32'd8030},
{32'd18132, -32'd3353, 32'd1932, -32'd14402},
{-32'd6520, -32'd8073, -32'd4677, -32'd968},
{-32'd5995, -32'd872, 32'd456, -32'd2011},
{32'd12404, 32'd5801, 32'd3486, 32'd3712},
{-32'd4304, -32'd4399, -32'd6694, -32'd74},
{-32'd1724, 32'd8171, -32'd5065, 32'd5469},
{32'd9895, -32'd844, -32'd4089, 32'd1951},
{-32'd10565, -32'd611, -32'd23234, -32'd2341},
{-32'd1480, -32'd1752, 32'd6955, 32'd1461},
{-32'd6003, -32'd1672, -32'd6357, -32'd4625},
{32'd1359, -32'd3746, -32'd749, -32'd9605},
{32'd2171, 32'd2109, -32'd6305, 32'd1519},
{-32'd11848, -32'd1210, -32'd5808, -32'd8471},
{-32'd12894, -32'd981, -32'd12071, -32'd4423},
{32'd1874, -32'd88, 32'd3471, -32'd3423},
{32'd9291, 32'd3957, 32'd747, 32'd2920},
{-32'd4653, -32'd1159, -32'd5588, 32'd655},
{-32'd1978, 32'd35, -32'd5678, -32'd4235},
{32'd398, -32'd8140, 32'd4283, -32'd3909},
{32'd4318, 32'd9160, -32'd1482, 32'd6131},
{32'd7824, -32'd1474, 32'd7846, -32'd3912},
{32'd2718, -32'd3782, -32'd8437, -32'd2411},
{32'd9421, -32'd5505, -32'd846, -32'd4279},
{32'd2141, 32'd189, 32'd6379, 32'd1536},
{-32'd13576, -32'd5408, -32'd4844, -32'd3500},
{32'd6712, 32'd5012, 32'd4824, 32'd9803},
{32'd7051, -32'd2901, 32'd855, 32'd4064},
{-32'd1918, -32'd1338, -32'd10778, -32'd3579},
{-32'd6663, 32'd2194, 32'd1381, -32'd106},
{32'd3996, 32'd8004, -32'd5713, -32'd5476},
{32'd1095, 32'd7347, -32'd18374, -32'd10164},
{-32'd3627, -32'd8443, -32'd4414, -32'd3584},
{-32'd12918, 32'd6033, -32'd13035, -32'd5578},
{-32'd3716, 32'd2060, 32'd6143, -32'd3809},
{32'd5153, -32'd534, 32'd9932, -32'd4075},
{32'd11028, 32'd2987, 32'd1202, 32'd4236},
{-32'd237, 32'd469, -32'd8216, -32'd5731},
{32'd10755, 32'd8745, 32'd11226, 32'd9269},
{-32'd5556, 32'd4546, -32'd3427, -32'd11371},
{-32'd4487, -32'd15070, -32'd4031, 32'd3591},
{-32'd7298, 32'd3183, 32'd9744, 32'd3769},
{32'd14649, 32'd15174, 32'd7310, 32'd842},
{32'd661, -32'd3654, -32'd5530, -32'd4342},
{-32'd3684, -32'd4612, -32'd10152, -32'd5532},
{32'd4944, -32'd8981, 32'd1070, 32'd653},
{32'd326, 32'd3057, 32'd3667, -32'd10737},
{-32'd125, -32'd5798, 32'd5020, -32'd10369},
{-32'd4803, 32'd2092, -32'd2811, 32'd6499},
{32'd12736, 32'd4082, 32'd3062, -32'd9993},
{-32'd1560, 32'd6021, 32'd4842, -32'd11594},
{32'd10534, 32'd6049, 32'd12562, 32'd7490},
{32'd2195, -32'd4331, 32'd7220, 32'd5279},
{-32'd4727, 32'd1451, 32'd1670, -32'd971},
{32'd10724, 32'd2203, 32'd6996, 32'd12545},
{32'd903, 32'd14651, 32'd4760, 32'd547},
{-32'd2713, -32'd3226, -32'd2715, 32'd9375},
{-32'd3511, -32'd7708, 32'd5051, -32'd2746},
{32'd2676, 32'd3133, 32'd11742, -32'd4004},
{32'd517, 32'd1898, -32'd8629, -32'd4768},
{-32'd16342, -32'd4776, -32'd8060, -32'd3411},
{-32'd2680, 32'd6008, -32'd4888, 32'd3943},
{32'd5142, 32'd187, -32'd3154, 32'd7505},
{32'd8523, -32'd200, 32'd1513, -32'd5622},
{-32'd9266, 32'd12030, -32'd3158, 32'd8231},
{-32'd6411, -32'd2238, -32'd7669, -32'd5526},
{32'd312, -32'd3119, -32'd7190, -32'd577},
{-32'd305, -32'd9136, -32'd23786, -32'd9598},
{-32'd3833, 32'd642, -32'd5542, -32'd3497},
{-32'd6829, -32'd6090, 32'd4183, -32'd1612},
{32'd7297, -32'd7124, 32'd2497, 32'd4687},
{-32'd1354, -32'd4684, 32'd484, -32'd7759},
{32'd5634, 32'd2710, 32'd7946, 32'd4664},
{-32'd1205, -32'd11278, -32'd15491, -32'd15269},
{32'd3529, 32'd13530, 32'd7305, 32'd2665},
{32'd14249, -32'd1346, 32'd14134, -32'd16503},
{-32'd868, -32'd841, -32'd6546, -32'd5643},
{32'd11546, -32'd10213, -32'd6355, 32'd2202},
{32'd4883, 32'd10492, -32'd6994, -32'd2901},
{32'd8055, -32'd2119, 32'd8143, 32'd11122},
{32'd4695, 32'd6089, 32'd7032, 32'd546},
{32'd1260, 32'd2246, -32'd3655, -32'd6352},
{32'd8091, 32'd10653, 32'd1496, 32'd597},
{32'd3613, -32'd6878, -32'd19902, 32'd430},
{-32'd5048, 32'd4104, 32'd2503, -32'd3401},
{-32'd4675, -32'd6417, -32'd7007, -32'd16207},
{32'd3631, 32'd3219, -32'd7736, -32'd13117},
{-32'd7814, 32'd1924, -32'd7573, -32'd7110},
{-32'd1358, -32'd1280, -32'd1850, 32'd3657},
{32'd11394, 32'd4787, -32'd2017, 32'd7646},
{32'd5175, 32'd8794, -32'd6926, 32'd5500},
{-32'd11118, -32'd261, 32'd1443, -32'd2111},
{-32'd9433, -32'd6604, -32'd1829, 32'd5158},
{-32'd8504, 32'd2551, -32'd488, -32'd6295},
{-32'd3801, -32'd5157, 32'd426, 32'd13103},
{-32'd647, 32'd2631, 32'd7912, -32'd5850},
{32'd8435, -32'd221, 32'd5302, 32'd1995},
{32'd2644, 32'd5099, -32'd6425, -32'd881}
},
{{32'd8781, 32'd5213, -32'd1712, -32'd2879},
{-32'd7741, -32'd12791, 32'd1163, -32'd18870},
{-32'd3564, 32'd4189, 32'd5025, -32'd6458},
{-32'd8308, -32'd3680, 32'd6695, 32'd9389},
{32'd221, 32'd491, 32'd3775, 32'd4888},
{32'd4117, -32'd5579, 32'd11570, 32'd8991},
{-32'd2347, 32'd4518, -32'd2704, -32'd1688},
{-32'd15222, 32'd7476, -32'd10487, -32'd1848},
{-32'd5516, 32'd7819, -32'd12865, -32'd11924},
{32'd3190, 32'd4902, -32'd39, -32'd4076},
{32'd4923, -32'd2077, 32'd7381, 32'd18894},
{32'd9090, 32'd3135, -32'd6065, 32'd5247},
{-32'd7647, -32'd1619, 32'd3690, 32'd8168},
{-32'd7306, -32'd4892, -32'd7303, 32'd1214},
{32'd5586, -32'd6723, -32'd6184, -32'd3036},
{32'd7226, -32'd9723, -32'd1825, 32'd13847},
{32'd512, 32'd17713, -32'd9559, 32'd2156},
{-32'd982, 32'd1788, 32'd3662, -32'd10694},
{-32'd21444, -32'd2753, -32'd1241, 32'd2487},
{32'd1821, -32'd13, 32'd109, -32'd6550},
{32'd1959, 32'd3567, -32'd2925, -32'd6536},
{-32'd7524, -32'd3952, 32'd9097, -32'd7928},
{32'd9916, 32'd5895, -32'd8439, -32'd5948},
{-32'd5348, -32'd6049, 32'd10373, 32'd6039},
{32'd6406, 32'd12716, 32'd11437, 32'd1610},
{-32'd12058, -32'd1153, 32'd9605, -32'd4133},
{32'd13378, 32'd7311, 32'd268, -32'd2872},
{-32'd6349, 32'd6358, -32'd4593, -32'd16690},
{-32'd845, 32'd8027, 32'd16295, 32'd3568},
{-32'd2885, -32'd1601, 32'd4673, 32'd4216},
{-32'd10021, 32'd2417, 32'd1873, 32'd3310},
{-32'd4968, -32'd4983, 32'd592, -32'd2420},
{32'd1849, 32'd8168, 32'd518, 32'd12582},
{-32'd1683, -32'd13271, -32'd4527, 32'd5307},
{32'd2009, 32'd7009, -32'd5120, -32'd8783},
{-32'd4825, 32'd1564, 32'd6072, -32'd8089},
{-32'd20254, -32'd2338, 32'd8713, -32'd2629},
{32'd1860, 32'd9034, -32'd6057, -32'd12652},
{-32'd5911, -32'd6381, -32'd10090, 32'd8101},
{32'd12972, -32'd1335, 32'd12103, 32'd9856},
{32'd1262, -32'd5824, 32'd624, -32'd3542},
{32'd3216, 32'd2455, 32'd868, -32'd9685},
{32'd17315, 32'd6334, 32'd2169, -32'd6584},
{-32'd152, -32'd674, -32'd10776, 32'd12902},
{-32'd2120, -32'd12695, -32'd2094, -32'd4438},
{-32'd815, -32'd6164, -32'd11452, -32'd1268},
{32'd8098, -32'd3471, 32'd6679, -32'd4454},
{32'd4651, -32'd14239, -32'd4784, 32'd17392},
{32'd1656, 32'd8015, 32'd7225, -32'd7629},
{-32'd1631, -32'd2898, -32'd8950, -32'd3302},
{32'd3816, -32'd4094, -32'd572, -32'd6360},
{32'd4657, 32'd2164, -32'd5018, 32'd1262},
{32'd6018, -32'd2226, -32'd1940, -32'd10740},
{32'd459, 32'd1454, 32'd16762, 32'd918},
{32'd5151, 32'd265, 32'd12825, 32'd13132},
{-32'd1580, 32'd3342, -32'd8392, -32'd16206},
{32'd111, 32'd5849, -32'd17623, 32'd20810},
{-32'd6791, -32'd15620, 32'd8001, 32'd5157},
{-32'd2417, -32'd3079, -32'd6025, -32'd5193},
{32'd176, 32'd5265, -32'd596, -32'd8994},
{-32'd9290, -32'd9349, 32'd1633, -32'd7332},
{-32'd12437, 32'd5475, -32'd3945, 32'd9004},
{-32'd6540, -32'd6279, -32'd1285, -32'd7116},
{-32'd7569, -32'd6091, -32'd206, -32'd8757},
{32'd47, -32'd184, -32'd1305, 32'd4083},
{32'd4479, 32'd4108, -32'd2319, 32'd3213},
{32'd8846, -32'd1191, -32'd8807, 32'd4841},
{32'd6639, 32'd1014, -32'd7572, -32'd5121},
{32'd8606, -32'd1074, -32'd9896, -32'd436},
{-32'd4609, 32'd3111, -32'd1769, -32'd14398},
{32'd1806, -32'd1711, 32'd4633, -32'd12222},
{-32'd8473, 32'd1071, 32'd15393, -32'd4872},
{32'd4471, -32'd3816, -32'd2177, -32'd3844},
{-32'd5628, -32'd2707, 32'd5989, 32'd1616},
{-32'd37, 32'd1341, 32'd4237, 32'd374},
{32'd15623, 32'd5752, -32'd2637, -32'd10894},
{-32'd10255, -32'd10090, 32'd2876, 32'd12443},
{-32'd3495, -32'd3437, -32'd10652, -32'd1544},
{-32'd3780, 32'd7696, 32'd7776, 32'd11329},
{32'd2225, 32'd13284, 32'd2243, -32'd2895},
{32'd279, -32'd4251, -32'd2052, 32'd16425},
{-32'd19799, 32'd238, 32'd1806, -32'd2614},
{-32'd15511, 32'd3530, 32'd5163, 32'd8626},
{32'd7965, 32'd5711, -32'd4660, 32'd2133},
{32'd14303, 32'd7101, 32'd6689, -32'd3616},
{32'd5133, -32'd4495, 32'd2599, -32'd5781},
{-32'd9277, -32'd2306, 32'd8116, 32'd1563},
{-32'd8648, -32'd4128, -32'd5915, 32'd1200},
{-32'd10428, -32'd2923, -32'd2449, 32'd7929},
{32'd2743, -32'd3958, 32'd8696, -32'd1883},
{32'd1674, 32'd10711, 32'd11890, 32'd12107},
{-32'd2877, -32'd14907, -32'd6955, -32'd7575},
{32'd4010, -32'd2246, 32'd15128, 32'd4166},
{32'd4761, -32'd1436, -32'd2324, 32'd673},
{32'd1420, 32'd6887, 32'd10901, 32'd1639},
{-32'd8165, 32'd3214, -32'd331, -32'd952},
{32'd541, 32'd4757, -32'd4227, 32'd3729},
{32'd15505, -32'd1998, 32'd22360, 32'd5710},
{-32'd8532, 32'd1574, 32'd16820, -32'd4762},
{32'd5737, 32'd3890, 32'd4151, -32'd8955},
{32'd8240, -32'd10748, 32'd1901, -32'd7936},
{-32'd231, -32'd7734, 32'd3451, -32'd13456},
{32'd266, 32'd6210, -32'd552, 32'd4707},
{32'd13356, 32'd4801, -32'd4990, 32'd4151},
{-32'd2726, 32'd890, -32'd530, 32'd2808},
{32'd2578, -32'd4122, -32'd7901, -32'd375},
{-32'd2511, -32'd2394, 32'd76, -32'd1359},
{32'd17899, 32'd921, -32'd13128, -32'd1856},
{32'd11137, 32'd4576, -32'd1775, 32'd2761},
{32'd3495, -32'd4772, 32'd10866, -32'd9775},
{-32'd3585, -32'd9527, -32'd5337, -32'd8219},
{32'd8529, 32'd10146, -32'd40, -32'd5513},
{32'd4844, 32'd6537, -32'd1782, 32'd13003},
{32'd2667, 32'd7175, -32'd7114, -32'd3478},
{32'd12336, -32'd9090, -32'd11579, -32'd2679},
{32'd2206, 32'd4629, -32'd5303, -32'd17162},
{32'd17386, 32'd7507, 32'd15170, -32'd4897},
{32'd8334, 32'd13612, 32'd2446, -32'd1855},
{-32'd13076, -32'd9461, -32'd5335, 32'd9735},
{-32'd1895, -32'd6399, -32'd3451, -32'd12094},
{32'd4878, 32'd7704, 32'd6595, 32'd254},
{-32'd10169, 32'd877, 32'd3611, 32'd4218},
{32'd15397, 32'd253, -32'd5568, 32'd665},
{-32'd10633, 32'd3409, 32'd7767, -32'd6540},
{-32'd3445, -32'd13460, 32'd8081, 32'd10668},
{32'd1885, 32'd5348, 32'd6666, -32'd5710},
{32'd4878, 32'd3255, -32'd8119, -32'd10585},
{-32'd10464, 32'd1001, -32'd4538, -32'd13841},
{32'd6098, -32'd9537, 32'd3734, -32'd6932},
{-32'd7129, 32'd11816, 32'd6453, -32'd10028},
{32'd3137, -32'd6400, -32'd1471, -32'd3216},
{32'd8755, -32'd8554, 32'd4992, 32'd6178},
{-32'd6886, -32'd13740, -32'd617, 32'd10997},
{-32'd3191, -32'd4561, 32'd6226, -32'd4663},
{-32'd587, 32'd1897, -32'd14660, 32'd4795},
{32'd2824, 32'd6243, -32'd11086, 32'd3463},
{-32'd3845, -32'd12566, 32'd4080, -32'd5402},
{-32'd6368, -32'd14069, -32'd3184, 32'd3536},
{32'd3091, 32'd4100, 32'd12378, -32'd5109},
{32'd9512, 32'd698, -32'd1293, -32'd1367},
{-32'd11165, -32'd1977, 32'd1715, 32'd6186},
{-32'd14678, 32'd2045, 32'd17086, -32'd1847},
{-32'd4474, -32'd7903, -32'd15872, 32'd7114},
{-32'd5404, 32'd5128, 32'd3189, 32'd8394},
{32'd225, 32'd3126, 32'd2340, -32'd7801},
{-32'd3931, 32'd7310, -32'd7234, -32'd4594},
{-32'd6753, 32'd406, -32'd8464, 32'd3864},
{-32'd7690, -32'd1594, 32'd7473, 32'd5261},
{32'd1767, 32'd393, 32'd2870, -32'd5388},
{32'd6866, 32'd3173, 32'd3564, 32'd9436},
{32'd1160, 32'd2434, 32'd2256, 32'd12078},
{-32'd5752, 32'd14269, 32'd857, -32'd140},
{32'd3796, 32'd4046, -32'd5474, -32'd4475},
{32'd658, -32'd2467, 32'd6500, 32'd6868},
{32'd642, 32'd2756, -32'd120, -32'd2784},
{32'd2493, -32'd8392, 32'd4748, 32'd2686},
{-32'd5746, 32'd1025, 32'd554, -32'd3614},
{-32'd2911, 32'd5412, -32'd15541, -32'd80},
{32'd7772, -32'd5603, -32'd3678, -32'd10092},
{-32'd5733, -32'd950, 32'd8373, 32'd3488},
{-32'd16728, 32'd6510, -32'd13166, 32'd2603},
{32'd156, 32'd16784, 32'd6612, -32'd257},
{-32'd7994, -32'd539, -32'd3706, -32'd19705},
{-32'd4954, 32'd8075, 32'd4732, 32'd6028},
{32'd10154, -32'd19025, 32'd20189, -32'd9140},
{-32'd4382, -32'd1144, -32'd10106, 32'd8075},
{32'd2535, -32'd2990, -32'd2278, 32'd3094},
{32'd2743, -32'd2645, 32'd8449, -32'd1831},
{32'd1133, -32'd12162, -32'd10678, 32'd8906},
{32'd5650, -32'd4464, 32'd2485, 32'd10979},
{-32'd6162, -32'd2787, -32'd3902, 32'd13089},
{32'd229, -32'd6611, 32'd13620, 32'd2060},
{32'd1464, 32'd1183, 32'd794, -32'd3734},
{-32'd5951, 32'd2666, 32'd8111, 32'd4928},
{32'd7905, 32'd3295, 32'd7265, -32'd13278},
{-32'd3569, -32'd2557, -32'd14177, 32'd857},
{-32'd223, 32'd4079, -32'd2104, 32'd2197},
{-32'd1897, 32'd11791, -32'd5052, -32'd3826},
{32'd11727, 32'd5245, 32'd9883, 32'd677},
{-32'd1528, -32'd15002, 32'd2341, 32'd13243},
{32'd1713, -32'd5096, -32'd1537, -32'd648},
{-32'd3970, 32'd882, 32'd1054, 32'd16358},
{32'd1824, 32'd1384, -32'd7597, 32'd15343},
{32'd5777, -32'd565, -32'd1340, 32'd281},
{32'd4442, 32'd1864, 32'd8104, 32'd222},
{32'd950, 32'd12217, -32'd5316, 32'd8679},
{-32'd1200, 32'd9497, 32'd9031, -32'd7355},
{32'd20815, 32'd14120, 32'd10719, 32'd2273},
{-32'd3311, -32'd427, -32'd920, 32'd9148},
{-32'd8879, 32'd1522, 32'd8495, 32'd2120},
{32'd10109, 32'd848, 32'd15341, 32'd3270},
{-32'd4784, -32'd13522, 32'd1592, 32'd2556},
{32'd21934, -32'd5622, 32'd4869, -32'd3270},
{-32'd1835, 32'd1921, 32'd17976, -32'd4154},
{32'd2255, -32'd1549, -32'd1046, -32'd13947},
{32'd17328, 32'd6809, -32'd151, -32'd5443},
{32'd7960, 32'd2015, -32'd14928, 32'd1265},
{32'd1982, -32'd1567, -32'd3518, -32'd1377},
{-32'd10178, -32'd8893, -32'd4776, 32'd4333},
{32'd4260, 32'd7685, -32'd12717, -32'd8714},
{-32'd5603, -32'd6245, 32'd4117, 32'd8639},
{32'd5850, -32'd1616, 32'd9518, -32'd2372},
{-32'd3888, 32'd2049, 32'd2329, 32'd4581},
{-32'd5143, 32'd4022, -32'd4664, 32'd2308},
{32'd5807, -32'd5315, 32'd2407, -32'd6788},
{-32'd12296, -32'd4656, 32'd6052, -32'd4790},
{32'd3810, -32'd5101, 32'd2892, -32'd1791},
{32'd7381, -32'd3229, -32'd6834, 32'd7812},
{-32'd6399, 32'd4627, -32'd10058, -32'd3355},
{32'd17682, 32'd2865, 32'd94, -32'd7834},
{32'd2456, -32'd4286, -32'd6037, -32'd10975},
{-32'd1184, -32'd3737, -32'd16078, -32'd15906},
{32'd1205, -32'd1451, 32'd5194, -32'd16309},
{32'd6514, -32'd2372, -32'd8035, -32'd8450},
{-32'd4098, -32'd3220, 32'd2561, -32'd1332},
{32'd9824, -32'd10063, -32'd3474, 32'd615},
{-32'd10933, -32'd1542, -32'd8824, -32'd11828},
{32'd1139, -32'd3648, -32'd10088, 32'd6278},
{-32'd6528, 32'd3713, 32'd8905, 32'd2115},
{32'd4515, -32'd93, -32'd7562, 32'd7606},
{32'd2845, -32'd8547, -32'd3562, 32'd4115},
{32'd313, 32'd8416, 32'd3865, -32'd1685},
{-32'd11696, 32'd514, 32'd5209, 32'd913},
{32'd86, 32'd1315, 32'd1538, 32'd7331},
{32'd6297, -32'd9677, 32'd7892, 32'd1841},
{-32'd5548, -32'd6049, -32'd3133, 32'd194},
{32'd1533, 32'd18277, -32'd1737, 32'd4995},
{-32'd5585, -32'd5567, -32'd9342, -32'd17666},
{32'd2904, -32'd2322, 32'd10275, -32'd4664},
{-32'd3604, 32'd2131, 32'd13550, 32'd3135},
{32'd4127, -32'd9352, -32'd9123, -32'd4778},
{32'd3438, -32'd1852, -32'd1180, -32'd10669},
{-32'd5600, -32'd3633, -32'd1872, -32'd1131},
{32'd7474, 32'd3172, 32'd7025, -32'd11064},
{-32'd1097, 32'd3725, 32'd1370, -32'd2737},
{-32'd8253, 32'd13328, 32'd5838, 32'd10256},
{32'd4172, -32'd6537, -32'd1597, -32'd6310},
{-32'd2487, -32'd9750, -32'd3693, 32'd8226},
{-32'd265, 32'd3505, 32'd3303, 32'd7530},
{32'd1772, -32'd3966, -32'd1138, 32'd694},
{32'd3757, -32'd10839, 32'd7909, -32'd716},
{-32'd5606, -32'd4932, -32'd10566, -32'd12551},
{-32'd7920, -32'd1496, 32'd6752, 32'd8570},
{32'd502, -32'd7790, 32'd1818, 32'd11418},
{32'd4447, 32'd392, -32'd7366, -32'd4390},
{-32'd3011, -32'd11739, -32'd6984, 32'd10741},
{32'd937, 32'd745, 32'd2157, 32'd1326},
{32'd7419, 32'd12598, 32'd6762, -32'd10822},
{32'd558, -32'd2355, -32'd1768, -32'd3536},
{32'd2695, 32'd13897, 32'd5269, -32'd1251},
{-32'd4597, -32'd6342, -32'd16768, 32'd4560},
{32'd6134, 32'd736, 32'd4661, -32'd59},
{-32'd4417, 32'd6169, 32'd9663, -32'd139},
{-32'd5313, -32'd7445, -32'd15062, 32'd9847},
{32'd2722, -32'd3962, -32'd2378, 32'd7407},
{-32'd1303, 32'd3237, -32'd9634, -32'd3252},
{32'd10628, 32'd734, -32'd6152, 32'd17937},
{32'd5142, -32'd4155, 32'd5588, 32'd9805},
{-32'd4734, -32'd5502, 32'd5616, 32'd13010},
{-32'd4212, 32'd1941, 32'd1909, -32'd3979},
{32'd3709, 32'd12207, -32'd7548, -32'd1040},
{-32'd3454, -32'd9138, -32'd835, -32'd8488},
{32'd1843, 32'd1235, 32'd2910, -32'd2149},
{32'd5064, -32'd11127, -32'd7064, 32'd8264},
{-32'd2479, 32'd12367, -32'd18, -32'd3555},
{-32'd16317, 32'd2518, -32'd9412, -32'd5695},
{-32'd10681, -32'd7241, 32'd8836, 32'd11360},
{-32'd2915, 32'd2291, 32'd15649, -32'd11266},
{-32'd5039, -32'd1569, 32'd3452, 32'd2690},
{-32'd10314, 32'd6825, -32'd9495, -32'd3105},
{-32'd8712, -32'd1486, -32'd14482, -32'd789},
{32'd3770, 32'd5079, -32'd4501, 32'd2586},
{-32'd2200, 32'd7666, -32'd5034, 32'd2051},
{32'd2177, 32'd1082, 32'd3989, -32'd10812},
{-32'd3482, -32'd937, -32'd15202, 32'd14342},
{-32'd13279, 32'd6461, 32'd2455, -32'd6217},
{32'd4748, 32'd4210, 32'd3154, -32'd4878},
{32'd5782, 32'd5040, -32'd1846, -32'd7452},
{32'd4671, 32'd4871, -32'd9260, 32'd3482},
{32'd8475, -32'd7640, -32'd4259, 32'd159},
{-32'd9222, 32'd8377, 32'd7247, 32'd91},
{-32'd1634, 32'd5310, 32'd522, -32'd11952},
{-32'd9570, 32'd10873, -32'd3299, 32'd10237},
{-32'd5421, -32'd14976, 32'd1279, 32'd5748},
{32'd7500, 32'd7280, 32'd4346, -32'd10451},
{-32'd12617, 32'd4802, 32'd637, 32'd11279},
{-32'd379, -32'd6130, 32'd4182, -32'd9331},
{32'd7280, 32'd3088, 32'd5238, 32'd5047},
{-32'd1490, 32'd5836, 32'd3857, -32'd7839},
{32'd8672, -32'd2645, -32'd443, 32'd2266},
{-32'd8824, -32'd17826, 32'd13375, 32'd10453},
{32'd5252, 32'd10240, 32'd8996, 32'd2618},
{-32'd89, -32'd1193, -32'd2641, -32'd6549},
{32'd10693, -32'd3586, 32'd2103, -32'd6994},
{32'd11006, -32'd8937, -32'd5856, 32'd1621},
{32'd8320, 32'd437, 32'd2783, 32'd9460},
{32'd11911, -32'd3058, 32'd3715, 32'd8959},
{32'd7931, 32'd7504, 32'd1611, -32'd14016},
{32'd7097, 32'd785, 32'd5570, 32'd2149},
{-32'd14392, 32'd1226, 32'd510, -32'd3312}
},
{{32'd8110, -32'd759, -32'd1515, 32'd483},
{-32'd3867, -32'd2149, 32'd4370, 32'd415},
{32'd7115, -32'd3259, 32'd4432, -32'd3187},
{-32'd6954, 32'd3043, 32'd9681, 32'd3925},
{-32'd2426, -32'd10663, -32'd4698, 32'd1253},
{-32'd5427, -32'd5483, 32'd1488, -32'd3706},
{-32'd9414, 32'd2205, -32'd5217, -32'd609},
{-32'd8291, -32'd577, -32'd5568, -32'd4589},
{-32'd6032, 32'd564, -32'd1143, 32'd634},
{32'd2813, 32'd5758, 32'd1745, 32'd5232},
{32'd9675, 32'd4372, -32'd3113, -32'd4046},
{-32'd373, 32'd4374, 32'd7934, -32'd3858},
{32'd5113, 32'd11707, -32'd2590, 32'd2392},
{32'd191, -32'd567, -32'd2136, 32'd2166},
{32'd1305, -32'd6032, -32'd1973, -32'd3806},
{32'd1717, -32'd11554, -32'd4740, -32'd899},
{32'd5607, -32'd6815, -32'd7348, 32'd6572},
{32'd1450, -32'd34, -32'd7217, -32'd350},
{-32'd12987, -32'd11442, -32'd2064, -32'd1780},
{-32'd9261, 32'd2631, -32'd6675, 32'd4},
{-32'd8509, 32'd14226, 32'd7519, -32'd1344},
{-32'd6486, -32'd6225, -32'd1309, -32'd2017},
{-32'd11243, -32'd1271, -32'd10140, 32'd4034},
{32'd4540, -32'd4048, -32'd4281, -32'd3511},
{32'd19015, 32'd7132, 32'd3930, 32'd270},
{32'd17687, -32'd190, 32'd3852, -32'd375},
{32'd7660, 32'd11201, 32'd2082, -32'd1768},
{-32'd3768, 32'd11246, -32'd9184, -32'd2115},
{32'd13828, -32'd1581, 32'd1548, 32'd5054},
{-32'd1523, -32'd1418, 32'd967, 32'd4074},
{32'd5996, -32'd3509, -32'd5701, 32'd6370},
{-32'd12903, -32'd4951, -32'd4930, -32'd3855},
{-32'd4920, 32'd3594, 32'd13279, 32'd3203},
{-32'd6152, -32'd337, 32'd1994, 32'd2686},
{32'd2310, 32'd1174, 32'd2739, 32'd6703},
{32'd14255, -32'd8772, -32'd10761, -32'd4058},
{32'd4800, -32'd7342, -32'd1312, 32'd1538},
{-32'd10610, -32'd13255, 32'd1940, 32'd6666},
{32'd2374, 32'd5457, -32'd294, 32'd2004},
{-32'd7151, -32'd3451, -32'd4451, -32'd2802},
{32'd10494, 32'd4155, -32'd534, 32'd1421},
{-32'd4835, 32'd8385, -32'd7726, 32'd800},
{32'd3475, -32'd1582, -32'd9118, -32'd1797},
{32'd1309, 32'd9992, -32'd1909, 32'd1116},
{-32'd10098, -32'd5656, -32'd6950, -32'd4356},
{32'd12103, 32'd2784, -32'd477, 32'd343},
{-32'd19297, -32'd3451, -32'd8759, -32'd3416},
{-32'd1468, -32'd12003, -32'd7120, 32'd4778},
{32'd3588, 32'd2366, -32'd935, 32'd5119},
{32'd5474, -32'd6480, -32'd453, 32'd2059},
{32'd415, 32'd7932, -32'd3546, 32'd339},
{32'd13759, 32'd12784, -32'd2243, 32'd1272},
{-32'd9568, 32'd5191, -32'd4125, 32'd196},
{-32'd5906, -32'd5580, -32'd7845, 32'd1650},
{32'd9342, 32'd488, -32'd4657, 32'd4493},
{-32'd7740, -32'd5463, 32'd10391, 32'd1855},
{-32'd4727, -32'd7359, -32'd2725, 32'd6091},
{-32'd10443, 32'd9459, 32'd2696, 32'd763},
{-32'd7685, -32'd6349, 32'd158, -32'd3010},
{-32'd10119, -32'd1436, -32'd1953, -32'd1710},
{32'd271, -32'd7584, -32'd195, -32'd1695},
{32'd2699, -32'd3570, 32'd694, -32'd2771},
{32'd2666, -32'd1768, -32'd6444, -32'd1473},
{32'd9674, 32'd6684, -32'd3632, 32'd1797},
{-32'd15700, -32'd1549, 32'd1876, -32'd1918},
{-32'd1366, 32'd13022, -32'd244, -32'd577},
{32'd1669, 32'd4032, 32'd10261, 32'd2660},
{-32'd12646, -32'd1401, -32'd561, -32'd2245},
{-32'd5799, -32'd2435, 32'd6399, -32'd2601},
{32'd2963, -32'd6691, 32'd3633, -32'd3258},
{32'd6117, 32'd1946, 32'd525, -32'd4844},
{32'd8490, -32'd5903, -32'd2229, -32'd1108},
{32'd4162, -32'd6842, -32'd2696, 32'd2168},
{-32'd15700, -32'd1121, 32'd1880, 32'd703},
{32'd6022, -32'd16, 32'd9028, 32'd6002},
{32'd25560, 32'd7617, -32'd9203, -32'd2058},
{32'd7586, 32'd94, -32'd669, 32'd2943},
{32'd6461, -32'd6517, 32'd3280, 32'd1592},
{32'd14051, 32'd4568, 32'd10799, 32'd1432},
{-32'd5876, 32'd4781, 32'd1261, 32'd5654},
{-32'd4307, -32'd5518, -32'd1506, -32'd102},
{-32'd13697, 32'd204, -32'd16196, -32'd1502},
{-32'd13744, -32'd10769, 32'd10087, -32'd1553},
{32'd513, 32'd8279, -32'd9478, 32'd5176},
{32'd4204, -32'd446, 32'd5767, -32'd3263},
{32'd71, -32'd8294, -32'd466, 32'd4170},
{32'd2729, -32'd6317, -32'd7230, -32'd1645},
{32'd1476, -32'd5706, -32'd15879, 32'd371},
{-32'd5535, 32'd47, 32'd8025, 32'd2184},
{-32'd11910, -32'd15758, 32'd2404, 32'd2016},
{32'd14005, -32'd5472, -32'd3072, -32'd1012},
{-32'd6566, 32'd3358, -32'd10448, 32'd3234},
{32'd3141, 32'd9638, -32'd4681, 32'd3524},
{32'd9811, 32'd11539, 32'd332, 32'd8046},
{32'd2527, 32'd3235, -32'd11073, 32'd6578},
{32'd8693, 32'd5513, -32'd10792, -32'd594},
{32'd48, -32'd835, 32'd1917, 32'd2245},
{32'd13541, -32'd5207, 32'd3957, 32'd6579},
{32'd980, 32'd4057, -32'd8226, 32'd1330},
{-32'd1349, 32'd6262, 32'd1954, -32'd948},
{32'd10104, -32'd1024, -32'd901, 32'd2142},
{32'd5284, -32'd6444, -32'd7790, 32'd940},
{-32'd7370, 32'd2602, -32'd88, 32'd1556},
{32'd9375, 32'd3350, 32'd7150, 32'd2935},
{32'd4880, -32'd10874, 32'd908, 32'd4109},
{-32'd5178, -32'd6008, 32'd1062, 32'd2914},
{-32'd12717, -32'd1109, -32'd7516, -32'd830},
{32'd16673, -32'd3091, -32'd1415, 32'd1527},
{32'd4681, 32'd4999, 32'd1484, -32'd2506},
{-32'd2852, 32'd2612, -32'd7728, 32'd3262},
{-32'd3338, -32'd4477, -32'd3600, -32'd4433},
{32'd3244, -32'd320, -32'd4576, -32'd2185},
{-32'd12731, -32'd2299, -32'd2674, 32'd3471},
{32'd2580, 32'd9530, 32'd4906, -32'd4489},
{-32'd1092, -32'd6301, 32'd8331, 32'd364},
{32'd3149, 32'd1358, 32'd4126, 32'd1172},
{32'd19740, -32'd1383, 32'd4608, 32'd1757},
{32'd6722, -32'd4420, -32'd3265, 32'd315},
{-32'd16340, -32'd5108, -32'd135, -32'd6414},
{-32'd9587, 32'd30, -32'd3748, 32'd803},
{-32'd3342, 32'd11160, 32'd8104, 32'd754},
{32'd2789, 32'd2953, 32'd9279, 32'd2235},
{32'd777, 32'd4954, 32'd2295, -32'd979},
{-32'd5525, -32'd8623, 32'd2806, -32'd1079},
{-32'd11973, -32'd10588, -32'd997, -32'd1134},
{-32'd211, 32'd420, -32'd1788, 32'd6141},
{-32'd1191, -32'd6766, 32'd3585, -32'd6561},
{-32'd2139, 32'd5025, -32'd15255, -32'd2119},
{-32'd14156, -32'd12406, -32'd10577, -32'd994},
{32'd6616, 32'd723, -32'd2912, -32'd231},
{-32'd4334, 32'd1344, -32'd7774, -32'd3581},
{-32'd11198, 32'd4273, 32'd6460, -32'd914},
{32'd5936, -32'd7249, -32'd4975, 32'd1778},
{32'd5981, 32'd2434, -32'd582, 32'd4237},
{-32'd5910, 32'd9419, 32'd6515, -32'd388},
{-32'd14477, -32'd9865, -32'd9950, 32'd2015},
{-32'd4771, 32'd3815, -32'd421, 32'd2870},
{32'd7906, 32'd11289, 32'd459, -32'd2435},
{-32'd10577, 32'd6353, 32'd3792, 32'd1296},
{32'd5555, -32'd6607, -32'd1258, -32'd1443},
{32'd2817, -32'd6112, -32'd9593, 32'd1027},
{-32'd6045, -32'd11581, -32'd10758, -32'd6883},
{-32'd1743, 32'd6612, 32'd795, 32'd2196},
{-32'd11492, -32'd3024, -32'd6888, 32'd2650},
{32'd6437, 32'd4032, 32'd2205, -32'd643},
{32'd42, -32'd1834, -32'd4266, 32'd1495},
{-32'd11940, 32'd852, -32'd7025, 32'd1867},
{32'd3312, -32'd2100, -32'd3413, 32'd1771},
{32'd3838, 32'd4931, -32'd1161, 32'd975},
{-32'd8852, -32'd12549, -32'd3692, -32'd5833},
{32'd3909, 32'd6437, -32'd5058, 32'd1007},
{32'd2305, -32'd2603, 32'd4413, 32'd7931},
{32'd4184, 32'd9289, 32'd7735, -32'd159},
{32'd16034, -32'd4172, -32'd1562, 32'd740},
{-32'd6908, -32'd11011, -32'd1255, -32'd4597},
{-32'd15765, -32'd724, 32'd3167, -32'd451},
{-32'd9156, 32'd3846, -32'd9790, 32'd4512},
{-32'd2948, -32'd3056, -32'd4674, 32'd1647},
{-32'd7749, 32'd2687, -32'd6319, -32'd519},
{-32'd3241, -32'd13599, 32'd2852, 32'd173},
{32'd5115, -32'd8907, -32'd3044, 32'd912},
{-32'd5940, 32'd12472, 32'd7854, -32'd785},
{32'd9543, -32'd4222, -32'd6493, -32'd2505},
{-32'd5245, 32'd4692, 32'd4995, -32'd4025},
{32'd17056, -32'd4417, -32'd742, 32'd4243},
{32'd2825, 32'd8877, 32'd664, 32'd1225},
{32'd7177, 32'd9237, 32'd4193, 32'd3820},
{32'd1822, -32'd4898, -32'd7098, -32'd4019},
{32'd3893, -32'd2405, -32'd1663, -32'd1111},
{-32'd5295, 32'd7984, 32'd2100, -32'd2348},
{-32'd17796, -32'd4980, 32'd6775, -32'd2277},
{-32'd6990, -32'd1415, 32'd2643, -32'd4142},
{-32'd5272, -32'd2400, -32'd2260, 32'd145},
{32'd4741, 32'd7659, -32'd2590, 32'd2011},
{-32'd376, -32'd14345, 32'd3100, -32'd1226},
{32'd1822, -32'd1461, 32'd8551, 32'd1929},
{32'd876, 32'd8442, 32'd2204, -32'd1702},
{32'd6651, -32'd8067, -32'd5984, 32'd6281},
{-32'd7520, -32'd8881, 32'd473, 32'd4269},
{-32'd12695, -32'd283, -32'd139, -32'd6895},
{-32'd5297, 32'd1824, -32'd6194, -32'd1949},
{-32'd13242, -32'd13592, -32'd10805, 32'd3997},
{-32'd2596, 32'd5657, -32'd558, -32'd7513},
{-32'd808, 32'd11046, 32'd1409, -32'd3135},
{-32'd10556, 32'd3665, -32'd6226, -32'd962},
{-32'd6926, 32'd3212, 32'd4872, 32'd3275},
{32'd3440, 32'd9079, -32'd1178, -32'd5272},
{-32'd10126, -32'd697, 32'd2973, -32'd1002},
{32'd3171, -32'd7335, -32'd11561, 32'd7652},
{-32'd648, -32'd1246, -32'd2462, -32'd2458},
{32'd5781, 32'd9062, 32'd1651, -32'd4180},
{-32'd2712, -32'd13217, -32'd4287, -32'd6697},
{-32'd16063, -32'd15198, -32'd16369, -32'd2301},
{32'd8349, -32'd1862, -32'd7465, 32'd4819},
{-32'd9677, 32'd111, 32'd244, -32'd941},
{32'd1316, -32'd7667, -32'd4953, -32'd2843},
{-32'd6422, -32'd1116, -32'd249, 32'd4760},
{-32'd1165, 32'd824, -32'd1396, 32'd651},
{-32'd17652, -32'd8096, 32'd9797, -32'd1419},
{-32'd4388, 32'd657, -32'd3416, -32'd3566},
{-32'd5643, -32'd10375, -32'd6503, -32'd1945},
{32'd648, 32'd6533, -32'd4189, -32'd3878},
{32'd9226, 32'd11538, -32'd97, -32'd4979},
{-32'd2902, 32'd8049, 32'd12348, 32'd2587},
{32'd1371, -32'd4358, 32'd2163, 32'd864},
{32'd6541, -32'd7868, -32'd2879, -32'd948},
{-32'd1595, 32'd3143, -32'd372, 32'd4956},
{-32'd2809, -32'd10787, -32'd2922, 32'd157},
{32'd1055, -32'd4509, 32'd8165, 32'd2412},
{32'd4272, -32'd9058, 32'd12503, 32'd1316},
{-32'd5688, -32'd4643, -32'd5356, 32'd2597},
{32'd58, 32'd10704, 32'd3336, 32'd4913},
{-32'd6119, -32'd7706, -32'd1445, -32'd4778},
{-32'd2115, 32'd8191, -32'd1415, -32'd5895},
{32'd16329, -32'd4918, -32'd1360, -32'd688},
{32'd8341, -32'd2780, 32'd155, -32'd1179},
{32'd1048, 32'd5302, 32'd5492, 32'd137},
{-32'd10312, 32'd10240, 32'd10497, -32'd1519},
{32'd9370, -32'd686, 32'd4456, 32'd3076},
{32'd687, 32'd15428, 32'd5741, -32'd2235},
{-32'd12035, 32'd2248, -32'd9088, 32'd2144},
{32'd14914, 32'd10736, 32'd7446, -32'd2136},
{-32'd3779, -32'd1496, 32'd1585, 32'd3919},
{32'd4383, 32'd9485, 32'd1845, -32'd8287},
{-32'd3961, 32'd3456, 32'd6498, -32'd2701},
{32'd3435, -32'd11123, 32'd4700, 32'd5575},
{-32'd15468, -32'd6821, -32'd1537, -32'd888},
{32'd11393, -32'd4356, -32'd14036, -32'd3858},
{-32'd15831, 32'd248, 32'd3281, -32'd1447},
{32'd13746, -32'd4051, 32'd1548, 32'd2148},
{32'd9224, -32'd4920, 32'd4616, -32'd1572},
{-32'd13078, 32'd2126, 32'd1869, -32'd3740},
{-32'd12222, -32'd681, 32'd175, -32'd178},
{32'd924, 32'd5618, 32'd2458, -32'd1238},
{-32'd6077, 32'd3666, 32'd4475, -32'd4713},
{32'd2431, 32'd4626, -32'd2654, -32'd4397},
{-32'd16536, -32'd8050, 32'd5495, 32'd4456},
{32'd4371, 32'd8728, 32'd1150, 32'd3848},
{-32'd6300, 32'd695, 32'd5416, -32'd2398},
{32'd5906, 32'd919, -32'd2789, 32'd1636},
{-32'd5081, -32'd151, 32'd1895, 32'd4043},
{32'd4072, -32'd1449, -32'd6347, 32'd2751},
{-32'd7186, -32'd2537, -32'd4399, -32'd6906},
{32'd13598, -32'd1567, -32'd425, 32'd5028},
{32'd4055, 32'd15765, 32'd8492, 32'd6236},
{32'd8579, 32'd5502, 32'd11670, -32'd2253},
{-32'd8947, -32'd6576, -32'd1330, -32'd3778},
{32'd5564, -32'd10834, -32'd7277, -32'd1010},
{-32'd4329, -32'd5717, 32'd3317, -32'd4240},
{32'd2887, 32'd2054, 32'd3725, 32'd4500},
{32'd4688, 32'd9490, 32'd7537, -32'd11},
{-32'd18358, -32'd2896, 32'd5387, 32'd1618},
{32'd14899, -32'd998, 32'd6988, 32'd3311},
{-32'd2074, 32'd296, 32'd3351, 32'd742},
{32'd5035, -32'd1272, -32'd2995, 32'd3904},
{-32'd2645, -32'd2804, -32'd3045, -32'd4784},
{-32'd9926, 32'd2540, 32'd622, 32'd3174},
{32'd10072, 32'd6029, 32'd9069, 32'd3317},
{-32'd7811, -32'd1584, -32'd4083, -32'd1270},
{-32'd2530, 32'd1041, 32'd10238, -32'd1144},
{-32'd6917, 32'd4254, 32'd6353, 32'd1428},
{-32'd2319, -32'd1440, 32'd6207, -32'd1982},
{32'd8679, -32'd12454, -32'd3489, -32'd5445},
{32'd1987, -32'd8297, -32'd2856, 32'd1037},
{-32'd6293, 32'd10098, 32'd377, 32'd558},
{-32'd6972, -32'd7726, 32'd834, 32'd617},
{32'd242, -32'd5430, 32'd3071, -32'd3418},
{32'd16988, -32'd1028, 32'd1431, -32'd156},
{-32'd8985, -32'd4808, -32'd12110, -32'd2886},
{32'd3367, -32'd7086, -32'd5235, 32'd4449},
{-32'd17789, -32'd4983, 32'd6748, 32'd2265},
{-32'd1394, 32'd2965, 32'd2225, 32'd3006},
{32'd17394, -32'd11181, -32'd9658, -32'd3602},
{32'd207, -32'd219, 32'd4693, 32'd1255},
{-32'd14951, 32'd3829, -32'd1013, 32'd4228},
{32'd8463, 32'd1191, -32'd7230, 32'd1667},
{32'd8233, 32'd9018, 32'd3192, 32'd1643},
{-32'd9153, 32'd8132, -32'd1088, -32'd2429},
{-32'd12146, -32'd10352, -32'd395, -32'd4045},
{-32'd251, -32'd12209, -32'd2262, -32'd496},
{-32'd9219, -32'd6446, 32'd577, 32'd1927},
{-32'd1885, 32'd12857, -32'd11398, 32'd3293},
{-32'd8173, -32'd2448, -32'd208, 32'd1849},
{-32'd13154, 32'd9304, 32'd1543, -32'd4193},
{32'd10015, -32'd265, -32'd8066, 32'd247},
{-32'd2911, -32'd7880, 32'd468, -32'd1167},
{-32'd1089, 32'd5855, 32'd5708, -32'd261},
{32'd195, 32'd2226, -32'd4603, -32'd2591},
{32'd3907, -32'd1507, -32'd9686, -32'd3271},
{32'd9840, 32'd467, 32'd3156, -32'd174},
{32'd10228, 32'd1052, -32'd3902, 32'd2691},
{32'd14227, 32'd3911, 32'd6537, -32'd2596},
{-32'd4476, -32'd3467, 32'd751, 32'd4604},
{32'd9263, -32'd1253, -32'd1805, -32'd4449},
{-32'd7735, -32'd4067, 32'd9132, -32'd7778},
{32'd1223, 32'd3531, 32'd2435, -32'd1685},
{-32'd1860, -32'd4293, -32'd4162, -32'd2606},
{32'd4138, 32'd8473, 32'd6262, -32'd16},
{-32'd377, 32'd4127, 32'd1506, -32'd2202},
{-32'd2671, -32'd7386, -32'd1957, -32'd3914}
},
{{-32'd2912, -32'd997, 32'd2115, -32'd10004},
{-32'd9180, 32'd286, -32'd16223, -32'd13051},
{-32'd7071, 32'd8483, -32'd10649, -32'd5242},
{32'd5859, -32'd6557, 32'd17748, -32'd297},
{-32'd606, -32'd6666, -32'd6663, -32'd14168},
{32'd3497, 32'd1682, -32'd4052, 32'd3476},
{32'd7371, 32'd6248, 32'd259, -32'd11175},
{-32'd9236, 32'd7216, -32'd2060, -32'd15379},
{-32'd7186, 32'd7022, -32'd6736, 32'd2789},
{32'd3403, 32'd1303, 32'd18334, 32'd9859},
{-32'd10065, -32'd1156, -32'd6171, 32'd5997},
{-32'd607, 32'd4212, 32'd1345, 32'd11442},
{-32'd272, -32'd7502, 32'd3702, 32'd17990},
{32'd18344, 32'd891, 32'd6988, -32'd740},
{-32'd5856, -32'd4532, 32'd6008, 32'd4917},
{-32'd3905, -32'd3331, 32'd1147, 32'd9339},
{32'd1461, -32'd5601, 32'd9068, 32'd4953},
{-32'd482, -32'd2968, -32'd7372, -32'd635},
{-32'd1721, 32'd8670, 32'd2912, -32'd3127},
{-32'd1041, -32'd8259, 32'd9185, -32'd12942},
{32'd11586, -32'd16906, -32'd4023, 32'd2477},
{32'd5707, 32'd1469, -32'd8059, -32'd10341},
{-32'd4333, -32'd8712, -32'd4388, 32'd6249},
{-32'd2358, 32'd7773, -32'd13645, -32'd12455},
{32'd2897, 32'd10528, 32'd16509, 32'd1098},
{32'd711, 32'd2678, -32'd12566, -32'd634},
{-32'd5120, -32'd14707, -32'd11872, 32'd4187},
{-32'd6313, 32'd7690, -32'd8826, 32'd2908},
{32'd393, 32'd3515, -32'd1112, -32'd6},
{32'd186, 32'd12827, -32'd6984, 32'd13294},
{32'd434, 32'd8431, 32'd5018, -32'd2374},
{-32'd3729, 32'd687, -32'd11424, -32'd9507},
{-32'd1395, -32'd7297, 32'd15254, -32'd90},
{-32'd3544, -32'd3979, -32'd4186, 32'd4633},
{32'd1930, 32'd2404, 32'd9561, 32'd3033},
{32'd602, 32'd3510, -32'd6488, -32'd15207},
{-32'd2491, 32'd4593, 32'd5335, -32'd3827},
{32'd50, -32'd7554, -32'd774, -32'd1185},
{-32'd11415, -32'd4716, 32'd3320, -32'd8343},
{-32'd4607, -32'd22027, 32'd6802, 32'd2017},
{-32'd1429, -32'd4048, -32'd300, -32'd1805},
{-32'd7389, -32'd3261, 32'd15802, 32'd9186},
{-32'd6452, -32'd3415, -32'd3056, -32'd15805},
{32'd4090, -32'd7713, 32'd2852, -32'd2134},
{32'd2853, 32'd1423, -32'd9419, -32'd10465},
{32'd3607, -32'd7160, 32'd6569, 32'd5167},
{32'd965, 32'd5323, -32'd13072, -32'd4070},
{-32'd10866, 32'd8791, -32'd940, -32'd2881},
{32'd8977, -32'd537, 32'd1428, 32'd3495},
{32'd5655, -32'd965, 32'd3904, -32'd3049},
{32'd3125, 32'd4155, -32'd10960, -32'd7623},
{-32'd949, -32'd6454, 32'd4457, 32'd1415},
{-32'd8286, -32'd4891, 32'd9460, -32'd15450},
{-32'd8346, 32'd6240, 32'd406, -32'd7258},
{32'd7540, -32'd5627, 32'd1318, -32'd4975},
{-32'd2117, 32'd7801, 32'd5838, 32'd1181},
{-32'd4773, -32'd9283, 32'd11473, 32'd3747},
{32'd4572, 32'd8108, -32'd20346, 32'd2239},
{-32'd6320, 32'd8829, -32'd13074, -32'd2797},
{-32'd10184, -32'd6690, -32'd8683, -32'd1282},
{-32'd8798, -32'd4499, -32'd14009, -32'd5901},
{-32'd17789, 32'd747, -32'd6092, 32'd13955},
{-32'd6652, -32'd3626, -32'd17874, -32'd14412},
{32'd1197, -32'd1845, -32'd1696, 32'd795},
{32'd13454, 32'd3926, 32'd15231, -32'd2865},
{-32'd3431, 32'd1910, 32'd2176, -32'd7728},
{32'd3468, -32'd3578, 32'd19042, 32'd9679},
{-32'd7361, -32'd6775, 32'd2513, -32'd4679},
{-32'd5720, 32'd5437, -32'd584, 32'd4799},
{32'd3451, 32'd5554, 32'd9377, -32'd916},
{-32'd2443, -32'd7732, 32'd6904, 32'd667},
{32'd8723, -32'd647, -32'd6417, -32'd9656},
{-32'd18734, -32'd4238, -32'd14952, 32'd6492},
{32'd314, -32'd4826, 32'd10234, -32'd19826},
{-32'd280, 32'd812, 32'd5071, -32'd1912},
{-32'd6193, -32'd2353, -32'd4387, 32'd13271},
{-32'd3717, 32'd4195, 32'd1250, -32'd7196},
{-32'd6544, 32'd3450, -32'd6722, 32'd8084},
{32'd1920, 32'd484, -32'd3048, 32'd3894},
{-32'd1262, -32'd10520, 32'd5511, -32'd5387},
{-32'd8625, -32'd13, -32'd2443, 32'd6018},
{-32'd1884, -32'd792, 32'd1268, -32'd4286},
{32'd10504, -32'd1925, -32'd10533, -32'd17078},
{32'd5010, -32'd1036, 32'd4137, -32'd3715},
{-32'd6668, 32'd5462, -32'd11070, -32'd3832},
{32'd6798, 32'd8379, 32'd11227, -32'd4335},
{-32'd190, 32'd3163, -32'd997, -32'd10131},
{-32'd1238, 32'd5144, -32'd12639, -32'd6989},
{-32'd3973, 32'd8626, 32'd1733, 32'd343},
{32'd1079, -32'd105, 32'd3249, -32'd9379},
{32'd4847, 32'd20, 32'd3963, 32'd341},
{-32'd2571, 32'd1935, -32'd7114, -32'd5378},
{-32'd7249, 32'd3190, -32'd6026, 32'd6212},
{-32'd5762, -32'd8585, 32'd9175, -32'd6754},
{32'd4116, 32'd11570, -32'd5688, -32'd6574},
{-32'd6142, 32'd9266, -32'd16097, -32'd10489},
{32'd672, -32'd380, 32'd1306, 32'd388},
{-32'd7738, 32'd861, 32'd10668, 32'd7728},
{32'd5388, 32'd10824, 32'd801, -32'd7304},
{-32'd3706, -32'd3306, 32'd3914, 32'd3579},
{-32'd3244, -32'd5126, 32'd13398, 32'd6997},
{32'd10385, 32'd10056, 32'd1262, -32'd3527},
{-32'd1997, 32'd412, 32'd1389, -32'd3407},
{-32'd1977, -32'd2346, 32'd3175, 32'd4759},
{32'd4684, -32'd6360, 32'd2373, 32'd5201},
{-32'd2050, 32'd3064, 32'd1103, -32'd3261},
{32'd5959, -32'd1898, -32'd5223, 32'd14278},
{32'd3924, -32'd6647, -32'd2340, 32'd3249},
{32'd16876, -32'd6454, 32'd3923, 32'd5945},
{-32'd8585, 32'd1439, -32'd5391, -32'd6814},
{-32'd8836, 32'd7357, -32'd10586, -32'd9980},
{-32'd9277, -32'd2817, 32'd1502, -32'd9917},
{32'd1397, -32'd14873, 32'd19054, 32'd3520},
{-32'd3352, -32'd13831, -32'd6088, 32'd1666},
{32'd3293, 32'd2711, -32'd5823, -32'd1011},
{-32'd2955, -32'd4168, -32'd4426, 32'd3186},
{32'd3807, 32'd9216, -32'd9895, 32'd2629},
{32'd1879, -32'd1032, -32'd8597, 32'd8804},
{32'd1112, 32'd1864, 32'd7756, -32'd15468},
{32'd481, -32'd5664, 32'd3610, 32'd4604},
{32'd6275, -32'd67, 32'd6919, -32'd16093},
{32'd423, 32'd4014, -32'd765, 32'd2337},
{-32'd3944, -32'd11384, -32'd6900, -32'd3592},
{32'd10254, 32'd14391, -32'd8149, -32'd9478},
{-32'd12280, -32'd7205, -32'd2273, -32'd8957},
{32'd5288, -32'd4235, 32'd9924, 32'd1672},
{-32'd4624, 32'd6836, -32'd9919, 32'd159},
{32'd133, 32'd8111, -32'd2777, -32'd9831},
{-32'd17428, 32'd8276, -32'd12457, 32'd4625},
{32'd1696, 32'd6800, -32'd15132, -32'd7580},
{32'd1319, 32'd6334, -32'd7930, -32'd7632},
{-32'd116, -32'd1132, -32'd8195, -32'd6887},
{32'd5237, -32'd677, -32'd4750, -32'd1158},
{32'd163, 32'd1972, -32'd4339, -32'd9185},
{32'd10507, 32'd7239, 32'd9837, 32'd12110},
{-32'd5985, 32'd6775, -32'd295, -32'd3540},
{32'd4281, 32'd12023, 32'd6933, 32'd6306},
{32'd4093, -32'd3105, 32'd3744, 32'd3362},
{-32'd2117, -32'd1717, 32'd10168, 32'd2703},
{32'd1093, -32'd9193, -32'd3863, -32'd6566},
{-32'd3002, -32'd5777, 32'd4878, -32'd7666},
{-32'd9061, 32'd4928, -32'd9032, 32'd2104},
{32'd3347, -32'd7639, -32'd8810, -32'd5095},
{-32'd579, 32'd11861, 32'd4073, 32'd3614},
{32'd1415, -32'd4451, 32'd3462, -32'd8944},
{-32'd5039, -32'd9587, 32'd5913, 32'd9341},
{-32'd681, -32'd15940, -32'd17013, -32'd1034},
{32'd6636, -32'd15124, 32'd9397, 32'd4276},
{-32'd4953, -32'd2286, 32'd6304, -32'd1117},
{-32'd6679, -32'd8198, -32'd8830, -32'd14831},
{32'd884, -32'd4372, -32'd3778, -32'd1012},
{32'd11748, -32'd3126, 32'd5406, -32'd6164},
{-32'd385, -32'd14713, -32'd2016, 32'd2892},
{-32'd8070, -32'd2544, 32'd3403, 32'd11326},
{32'd1283, 32'd3000, -32'd2455, -32'd688},
{32'd8022, 32'd5664, 32'd559, 32'd10942},
{32'd7062, 32'd2842, -32'd313, 32'd2969},
{32'd6539, 32'd8619, 32'd8018, 32'd6970},
{-32'd11210, -32'd10318, -32'd7907, -32'd9623},
{32'd1752, 32'd4006, -32'd2310, -32'd2102},
{-32'd3641, 32'd10587, -32'd10514, -32'd13375},
{32'd3266, -32'd2151, 32'd8005, -32'd828},
{32'd751, -32'd8089, -32'd5266, 32'd2294},
{-32'd2516, 32'd9048, 32'd11424, -32'd11418},
{32'd5176, -32'd1027, 32'd5214, 32'd3868},
{-32'd4401, -32'd11468, 32'd15831, 32'd1357},
{32'd17357, 32'd1292, 32'd1961, 32'd716},
{-32'd10127, 32'd6720, -32'd26690, -32'd4701},
{32'd4788, -32'd8044, -32'd18157, 32'd3209},
{-32'd3295, 32'd1760, -32'd11175, -32'd2462},
{-32'd6590, 32'd3051, 32'd2272, 32'd2898},
{32'd4680, -32'd1970, 32'd2840, -32'd8554},
{32'd12879, 32'd2054, 32'd9473, 32'd1591},
{-32'd14291, -32'd789, 32'd438, 32'd4900},
{32'd8046, 32'd2230, -32'd4136, -32'd8300},
{32'd15102, 32'd436, 32'd7268, 32'd422},
{32'd7207, -32'd295, 32'd7352, 32'd10496},
{32'd1366, -32'd4589, 32'd7937, 32'd6248},
{32'd6737, -32'd1434, -32'd787, -32'd8431},
{-32'd10372, -32'd5869, -32'd1262, 32'd1609},
{-32'd8293, -32'd6892, -32'd4445, 32'd868},
{32'd2655, -32'd6809, -32'd3437, -32'd1090},
{32'd1107, -32'd7246, 32'd9425, 32'd5500},
{-32'd11614, -32'd7241, -32'd2937, 32'd442},
{32'd12147, -32'd2083, -32'd1743, 32'd2578},
{32'd6365, -32'd1463, 32'd10217, 32'd8501},
{32'd3703, 32'd2338, -32'd4445, 32'd416},
{-32'd1293, -32'd3925, 32'd8391, 32'd3666},
{-32'd10287, 32'd224, -32'd7963, 32'd7516},
{32'd13304, 32'd7745, -32'd2466, 32'd9519},
{-32'd289, -32'd5904, 32'd10926, -32'd8500},
{32'd1653, -32'd709, -32'd3836, -32'd1294},
{32'd5577, -32'd5319, -32'd100, 32'd954},
{-32'd4135, -32'd431, 32'd2372, -32'd4741},
{32'd1138, 32'd2758, 32'd3464, -32'd5632},
{-32'd15692, -32'd13723, -32'd12820, -32'd1924},
{32'd2401, -32'd10502, -32'd4914, 32'd10987},
{-32'd2962, -32'd2277, 32'd4528, 32'd2665},
{-32'd8904, 32'd15157, -32'd8650, 32'd511},
{32'd1836, 32'd4391, 32'd7812, 32'd4532},
{32'd4934, 32'd1128, -32'd6245, 32'd1317},
{-32'd9213, -32'd197, -32'd2549, -32'd336},
{-32'd4196, -32'd2790, -32'd4844, -32'd11682},
{32'd459, -32'd6777, 32'd11135, -32'd10652},
{-32'd12131, 32'd3733, -32'd6831, 32'd9200},
{32'd9533, 32'd3985, -32'd5108, 32'd5977},
{32'd3381, 32'd2513, 32'd9069, 32'd7385},
{-32'd10465, -32'd2924, 32'd5148, -32'd7974},
{-32'd572, 32'd12667, -32'd13119, -32'd285},
{32'd6058, 32'd5800, -32'd5073, -32'd9192},
{-32'd15740, -32'd13305, 32'd285, -32'd5452},
{32'd6942, 32'd8, -32'd1697, -32'd5569},
{-32'd4426, 32'd9722, -32'd2962, -32'd18586},
{-32'd14010, -32'd7469, -32'd6896, 32'd11014},
{32'd726, -32'd14629, 32'd135, -32'd983},
{32'd5026, -32'd4597, 32'd4406, 32'd2648},
{32'd4591, 32'd5217, -32'd942, -32'd3393},
{32'd4584, 32'd1338, -32'd4306, -32'd3249},
{32'd13140, -32'd9526, 32'd9931, 32'd1277},
{-32'd5272, -32'd3401, -32'd3757, 32'd7111},
{-32'd431, 32'd3282, 32'd6125, 32'd12801},
{32'd2963, -32'd5262, 32'd3816, -32'd4799},
{-32'd6896, 32'd11324, -32'd425, 32'd3534},
{32'd397, 32'd15746, 32'd3592, 32'd10905},
{-32'd2760, -32'd1478, -32'd2373, -32'd1352},
{-32'd2354, -32'd6202, -32'd9142, -32'd19334},
{32'd736, 32'd9729, 32'd1491, 32'd5630},
{-32'd14208, 32'd9542, -32'd9048, -32'd14990},
{-32'd2070, 32'd7298, 32'd10655, 32'd2541},
{32'd13257, -32'd2164, 32'd15601, -32'd1494},
{-32'd2605, -32'd1973, -32'd14810, 32'd5259},
{-32'd7037, 32'd10845, 32'd4586, -32'd6765},
{-32'd15069, 32'd2759, -32'd2303, 32'd3282},
{-32'd7385, 32'd3003, -32'd3140, -32'd11812},
{32'd2790, -32'd6106, -32'd5024, 32'd6562},
{-32'd4046, 32'd1146, -32'd12332, 32'd2896},
{32'd5611, 32'd8090, 32'd5296, 32'd2322},
{-32'd4688, 32'd5251, -32'd7855, 32'd3738},
{32'd8632, 32'd3877, 32'd3535, 32'd14880},
{32'd2480, 32'd10704, -32'd14491, 32'd3625},
{32'd2473, -32'd10647, -32'd507, -32'd4650},
{-32'd5991, 32'd7016, 32'd5704, -32'd3021},
{-32'd2979, -32'd2624, -32'd13532, -32'd10340},
{32'd2909, 32'd1611, 32'd10014, 32'd5409},
{32'd2855, 32'd2849, 32'd17749, 32'd6983},
{-32'd3469, 32'd6214, -32'd849, -32'd10346},
{-32'd2106, 32'd6308, -32'd15454, -32'd10518},
{32'd1514, 32'd3221, 32'd2899, 32'd1051},
{-32'd3159, 32'd7692, -32'd8756, -32'd3877},
{-32'd3945, -32'd6538, -32'd9615, 32'd6880},
{-32'd7735, 32'd884, 32'd756, -32'd11181},
{32'd5043, 32'd5449, -32'd1346, 32'd6064},
{32'd17659, 32'd8673, 32'd7005, 32'd10429},
{-32'd5413, -32'd6740, 32'd17998, -32'd1821},
{-32'd423, 32'd971, -32'd5410, -32'd5944},
{32'd7395, 32'd4522, -32'd1400, -32'd3534},
{-32'd2450, -32'd4789, 32'd11909, -32'd1832},
{32'd847, -32'd777, 32'd19675, -32'd6312},
{-32'd4669, -32'd7254, -32'd3514, -32'd5306},
{32'd489, -32'd1091, -32'd1095, 32'd7124},
{32'd9182, 32'd3927, 32'd9628, 32'd1049},
{32'd15344, 32'd7869, 32'd1049, -32'd6019},
{-32'd1909, 32'd4855, -32'd6481, 32'd1003},
{-32'd6197, 32'd6121, -32'd1543, 32'd1569},
{-32'd5433, -32'd320, 32'd2034, -32'd2449},
{-32'd10143, 32'd6316, -32'd3727, 32'd547},
{32'd3999, -32'd57, 32'd6750, 32'd6790},
{32'd2398, -32'd5196, 32'd2381, -32'd6970},
{32'd2211, 32'd10503, -32'd7380, -32'd3454},
{32'd4002, -32'd5482, -32'd8400, -32'd10710},
{-32'd9539, 32'd4288, 32'd6387, -32'd107},
{32'd1160, 32'd3491, 32'd5765, -32'd8428},
{-32'd5039, 32'd1404, -32'd7060, -32'd2769},
{-32'd3660, -32'd1519, 32'd8269, 32'd16509},
{-32'd3584, 32'd4140, 32'd937, -32'd5098},
{-32'd10114, 32'd4024, -32'd8261, -32'd12772},
{32'd4193, 32'd2249, 32'd13650, 32'd3695},
{32'd1866, 32'd1862, -32'd18625, 32'd17995},
{-32'd1968, 32'd8985, -32'd10862, -32'd218},
{32'd7360, 32'd7035, 32'd4893, 32'd2928},
{-32'd2502, 32'd7614, 32'd7296, -32'd2200},
{32'd1933, 32'd4337, -32'd3988, -32'd1832},
{-32'd3193, 32'd7854, 32'd6338, 32'd8692},
{-32'd2974, -32'd1906, 32'd4963, -32'd65},
{-32'd2563, 32'd1703, -32'd4816, 32'd672},
{-32'd8946, -32'd3892, -32'd10956, -32'd6501},
{-32'd10514, 32'd3956, -32'd2321, -32'd4019},
{-32'd2383, -32'd3154, 32'd6934, 32'd8466},
{-32'd2380, 32'd15904, -32'd5810, -32'd11650},
{-32'd10907, 32'd5869, -32'd2240, -32'd19252},
{32'd4461, 32'd2206, -32'd5501, -32'd2065},
{-32'd4617, -32'd658, 32'd7317, -32'd2337},
{-32'd4456, 32'd4924, -32'd4238, 32'd1819},
{32'd1010, 32'd7920, -32'd15125, -32'd1391},
{32'd1595, 32'd2754, -32'd6353, 32'd1753},
{32'd4594, -32'd11517, 32'd2279, -32'd66},
{32'd10674, -32'd3189, 32'd1884, 32'd5672},
{32'd9540, 32'd1717, 32'd4993, 32'd9349},
{32'd3228, 32'd4816, 32'd11514, -32'd4608},
{32'd927, 32'd1455, -32'd4988, -32'd5279}
},
{{-32'd958, 32'd1458, 32'd1221, -32'd3454},
{-32'd1119, -32'd12297, 32'd10253, 32'd5715},
{32'd8484, -32'd1544, -32'd16711, -32'd6072},
{32'd9365, 32'd1793, 32'd215, -32'd7222},
{32'd8940, -32'd5895, 32'd4801, -32'd3164},
{32'd2445, -32'd4216, 32'd5008, -32'd3420},
{-32'd9614, -32'd1864, -32'd6793, -32'd6631},
{32'd7712, -32'd6427, 32'd1316, 32'd1428},
{32'd9319, 32'd11003, -32'd2520, 32'd5159},
{32'd4436, 32'd6796, -32'd8729, -32'd3526},
{32'd288, -32'd11509, -32'd4564, -32'd1509},
{-32'd2088, -32'd1589, 32'd12547, 32'd5457},
{-32'd622, -32'd3957, -32'd5049, -32'd12820},
{-32'd3726, -32'd5103, 32'd2238, -32'd950},
{-32'd7242, -32'd7564, 32'd2329, 32'd1478},
{-32'd485, 32'd2162, 32'd8167, -32'd6453},
{32'd2313, -32'd3393, 32'd14828, 32'd4311},
{32'd12182, 32'd8517, -32'd6935, 32'd3242},
{32'd10061, 32'd9212, -32'd5878, -32'd6601},
{-32'd1146, 32'd3235, -32'd348, 32'd5246},
{-32'd1935, 32'd1447, -32'd2640, -32'd1439},
{-32'd2692, -32'd5178, 32'd6093, 32'd3666},
{32'd11208, 32'd5821, 32'd8113, 32'd9615},
{32'd6871, 32'd4933, -32'd7751, -32'd1345},
{32'd421, 32'd3032, -32'd8184, -32'd4692},
{-32'd2479, -32'd7679, -32'd4396, -32'd153},
{-32'd1697, 32'd3821, 32'd14757, -32'd1649},
{32'd4544, 32'd12276, -32'd2526, -32'd2157},
{32'd10129, -32'd8231, 32'd5300, -32'd6643},
{-32'd10950, -32'd1954, -32'd17297, 32'd11146},
{-32'd5838, -32'd3618, 32'd10945, -32'd2587},
{-32'd3971, -32'd8545, 32'd9615, 32'd5637},
{-32'd405, -32'd2177, 32'd3472, 32'd575},
{32'd4578, 32'd6715, 32'd2201, 32'd3800},
{32'd749, 32'd1985, -32'd6819, -32'd7424},
{-32'd10409, -32'd19255, -32'd16685, -32'd4938},
{32'd1540, -32'd5140, -32'd836, -32'd3437},
{32'd3168, 32'd5089, 32'd1405, 32'd5984},
{32'd2633, 32'd2512, 32'd8057, -32'd10446},
{32'd3979, 32'd1118, -32'd10980, 32'd8623},
{32'd394, 32'd11378, -32'd8460, -32'd447},
{32'd1024, -32'd4209, -32'd13482, 32'd5040},
{32'd1167, 32'd1198, -32'd13170, 32'd6605},
{-32'd3374, 32'd190, 32'd6067, -32'd2676},
{-32'd1473, 32'd5583, -32'd480, 32'd3315},
{-32'd2907, 32'd6048, 32'd7481, -32'd429},
{-32'd12752, 32'd1537, -32'd9234, 32'd6296},
{32'd3695, 32'd4124, 32'd6843, 32'd13813},
{-32'd2492, -32'd4882, -32'd13427, -32'd768},
{-32'd1394, -32'd1994, 32'd6538, 32'd7279},
{-32'd4619, -32'd766, 32'd14423, 32'd8144},
{-32'd2839, -32'd10151, 32'd3347, -32'd3619},
{-32'd1403, 32'd3932, 32'd6696, 32'd8156},
{-32'd1727, -32'd4372, -32'd2832, 32'd6487},
{32'd4992, -32'd4434, 32'd1212, -32'd7119},
{32'd780, -32'd11135, 32'd8661, -32'd1600},
{-32'd960, 32'd6369, -32'd3726, -32'd2944},
{-32'd17989, 32'd1037, 32'd2536, -32'd1012},
{32'd4096, -32'd1498, 32'd7088, -32'd6893},
{-32'd1333, 32'd3242, 32'd2141, -32'd3153},
{32'd7438, -32'd7236, -32'd2841, 32'd741},
{32'd8351, 32'd3970, -32'd8972, 32'd3107},
{-32'd1613, -32'd2070, 32'd4324, -32'd86},
{-32'd10848, -32'd15984, 32'd7220, 32'd4284},
{32'd8866, 32'd8717, -32'd2611, 32'd7974},
{32'd6833, -32'd7463, 32'd1375, -32'd4200},
{-32'd3065, -32'd5593, 32'd19119, 32'd1348},
{32'd9934, 32'd1827, 32'd1090, 32'd9755},
{32'd8934, 32'd98, 32'd4329, 32'd7647},
{-32'd7131, -32'd2066, -32'd166, -32'd5719},
{-32'd10339, -32'd78, 32'd9941, -32'd9861},
{32'd4193, -32'd6252, 32'd1221, -32'd5105},
{-32'd11372, 32'd7628, 32'd7304, -32'd1669},
{32'd1205, -32'd10683, 32'd12291, 32'd16747},
{32'd12014, 32'd5569, 32'd3508, 32'd8300},
{32'd6438, 32'd6614, -32'd445, 32'd4873},
{32'd1674, -32'd596, 32'd4706, 32'd2155},
{-32'd4396, 32'd250, 32'd7470, 32'd3504},
{-32'd1587, 32'd1763, -32'd4088, -32'd11079},
{-32'd2646, -32'd6493, 32'd4699, -32'd9069},
{32'd11973, 32'd4617, -32'd2072, -32'd12591},
{-32'd8351, -32'd258, 32'd2747, -32'd5183},
{32'd4761, -32'd562, 32'd3960, -32'd7491},
{32'd10985, 32'd103, 32'd10699, 32'd4793},
{-32'd4141, -32'd5444, -32'd4451, 32'd2422},
{32'd8781, -32'd837, 32'd18318, 32'd1419},
{-32'd758, 32'd9508, -32'd11875, 32'd3620},
{-32'd5399, -32'd5110, 32'd11733, -32'd6968},
{32'd6127, 32'd4674, 32'd5242, -32'd1543},
{32'd2074, 32'd710, 32'd1121, 32'd1545},
{-32'd890, 32'd3475, -32'd16786, 32'd8551},
{32'd8245, -32'd396, -32'd2997, 32'd14432},
{32'd6662, 32'd4423, -32'd6975, 32'd861},
{32'd5144, -32'd1823, 32'd3458, 32'd690},
{32'd3890, -32'd1907, -32'd2854, 32'd6943},
{-32'd9981, 32'd1507, -32'd1630, -32'd4582},
{32'd7628, 32'd8839, -32'd7929, -32'd654},
{32'd6247, 32'd2221, -32'd5750, -32'd2835},
{-32'd713, -32'd4983, -32'd4345, 32'd15306},
{-32'd907, 32'd5055, -32'd6138, 32'd3129},
{-32'd16622, 32'd3066, -32'd1770, -32'd4256},
{32'd10252, 32'd2661, 32'd733, 32'd365},
{32'd1035, 32'd10512, -32'd1761, 32'd2092},
{32'd6287, 32'd16424, 32'd23183, 32'd890},
{-32'd882, 32'd1375, 32'd6816, 32'd5239},
{-32'd10551, 32'd4579, -32'd4441, 32'd1049},
{-32'd6381, -32'd1819, -32'd13610, -32'd2565},
{32'd5395, -32'd559, 32'd7032, 32'd2405},
{-32'd790, 32'd7731, -32'd612, -32'd6256},
{-32'd8788, -32'd3744, 32'd6100, 32'd7652},
{-32'd2423, 32'd9643, 32'd12060, -32'd2934},
{32'd1774, -32'd7917, 32'd4273, -32'd3326},
{32'd1914, 32'd374, 32'd3684, 32'd2197},
{32'd784, -32'd5068, -32'd7341, -32'd2554},
{-32'd4026, 32'd10470, 32'd1658, 32'd2253},
{32'd55, 32'd2534, 32'd13861, 32'd8583},
{32'd6493, 32'd2533, -32'd5085, 32'd7738},
{32'd2657, 32'd524, -32'd4909, 32'd6968},
{-32'd9425, -32'd8966, 32'd14607, -32'd12709},
{-32'd11475, -32'd927, -32'd2729, -32'd4151},
{32'd5226, 32'd3167, 32'd9120, 32'd2545},
{32'd3665, 32'd15780, -32'd3803, 32'd4751},
{32'd6622, -32'd13423, 32'd21478, -32'd2567},
{32'd6237, 32'd12805, -32'd783, 32'd2050},
{-32'd8865, -32'd6303, -32'd15213, 32'd8156},
{32'd715, 32'd2436, -32'd3033, 32'd11231},
{-32'd3425, 32'd5480, -32'd2826, 32'd5998},
{32'd7574, 32'd1107, 32'd4447, 32'd251},
{-32'd1216, 32'd9200, -32'd5431, 32'd13441},
{32'd1690, -32'd5810, 32'd1901, 32'd235},
{32'd3134, -32'd2871, 32'd12505, 32'd9304},
{32'd6185, 32'd1641, 32'd8343, 32'd10248},
{-32'd3497, 32'd7425, -32'd308, -32'd9143},
{-32'd5304, -32'd5435, -32'd1567, -32'd2672},
{32'd3451, 32'd18843, 32'd8720, -32'd1411},
{32'd703, -32'd5304, 32'd12633, -32'd4367},
{-32'd1689, 32'd5175, 32'd5368, -32'd5331},
{-32'd5780, 32'd8427, 32'd2122, -32'd6874},
{32'd9426, -32'd3816, -32'd5743, 32'd3123},
{-32'd1347, 32'd1856, 32'd1524, 32'd2220},
{-32'd6613, -32'd1266, 32'd10612, 32'd4014},
{32'd6353, -32'd12668, -32'd7694, -32'd11863},
{32'd4779, -32'd8001, 32'd5287, -32'd4181},
{-32'd7355, 32'd578, 32'd3941, 32'd3478},
{-32'd5067, -32'd4126, -32'd6113, -32'd8010},
{32'd5441, -32'd4160, 32'd491, 32'd6941},
{32'd12678, -32'd2554, -32'd5291, 32'd4090},
{-32'd7460, -32'd872, -32'd2614, -32'd5},
{-32'd8511, -32'd8156, -32'd7957, 32'd410},
{32'd1646, -32'd8538, 32'd7442, -32'd5157},
{32'd2081, 32'd2760, -32'd301, -32'd4281},
{32'd10794, 32'd1020, 32'd4384, -32'd6847},
{-32'd2444, -32'd1781, 32'd13574, 32'd7371},
{32'd6744, -32'd738, 32'd2806, -32'd2559},
{32'd4962, 32'd851, -32'd4637, 32'd8222},
{-32'd4980, 32'd19414, -32'd1839, 32'd2441},
{32'd5319, 32'd430, -32'd1617, -32'd3786},
{32'd14720, -32'd3162, -32'd6792, 32'd3811},
{32'd5912, 32'd4562, 32'd11468, 32'd5334},
{32'd942, -32'd5967, -32'd17309, 32'd6506},
{-32'd213, 32'd3192, 32'd18183, 32'd6273},
{32'd6403, 32'd6643, -32'd2910, -32'd9258},
{32'd2726, -32'd1429, 32'd3548, 32'd3555},
{-32'd2082, -32'd16018, -32'd3698, -32'd6891},
{32'd707, -32'd1911, -32'd12523, -32'd3346},
{-32'd728, 32'd1899, 32'd8060, 32'd1520},
{-32'd13319, 32'd3319, -32'd9173, 32'd10367},
{32'd7621, -32'd1244, 32'd13357, -32'd4929},
{-32'd11022, -32'd1918, -32'd5860, -32'd7650},
{-32'd2617, -32'd1241, 32'd1851, 32'd7948},
{-32'd10852, -32'd2982, -32'd6694, 32'd7273},
{-32'd17051, 32'd3050, -32'd12229, 32'd726},
{32'd6490, 32'd587, -32'd6120, -32'd3040},
{32'd3721, 32'd3400, -32'd8116, 32'd364},
{-32'd262, -32'd13284, -32'd2889, -32'd5348},
{32'd95, -32'd6747, -32'd1464, 32'd5398},
{32'd3030, 32'd14487, -32'd5597, -32'd1269},
{-32'd7269, -32'd2392, 32'd10595, -32'd7459},
{-32'd6606, 32'd2511, 32'd7944, 32'd579},
{-32'd4816, 32'd6295, 32'd1994, 32'd8223},
{32'd1147, -32'd4818, 32'd13411, 32'd5808},
{32'd797, 32'd1883, 32'd9527, 32'd1605},
{-32'd6792, -32'd2937, -32'd2345, -32'd2652},
{-32'd8206, 32'd11337, 32'd1422, 32'd4967},
{-32'd3432, -32'd8154, -32'd7909, -32'd8543},
{-32'd658, -32'd3204, -32'd103, 32'd2270},
{32'd824, -32'd13510, -32'd11331, -32'd2684},
{-32'd9385, 32'd488, 32'd17237, 32'd6757},
{-32'd2107, 32'd7871, 32'd13753, -32'd9689},
{32'd741, 32'd2278, 32'd2251, -32'd20021},
{-32'd2298, -32'd10067, -32'd9029, -32'd4291},
{-32'd10423, -32'd2538, 32'd5574, -32'd7815},
{-32'd1066, 32'd6050, -32'd1134, -32'd380},
{32'd924, 32'd4092, -32'd1682, -32'd11005},
{32'd2908, 32'd3914, 32'd11889, 32'd8597},
{-32'd670, 32'd3005, 32'd598, 32'd4829},
{-32'd11233, 32'd1392, 32'd10693, -32'd9630},
{32'd11398, -32'd4630, 32'd13693, -32'd5651},
{-32'd6431, 32'd4430, 32'd2469, -32'd236},
{-32'd3404, 32'd9258, -32'd5880, 32'd1726},
{-32'd854, 32'd1803, -32'd573, 32'd12844},
{-32'd6761, 32'd548, -32'd1163, 32'd5892},
{32'd10720, 32'd1725, 32'd3014, 32'd3044},
{32'd3162, -32'd4593, 32'd19136, -32'd6610},
{-32'd48, -32'd2344, 32'd8395, -32'd4138},
{-32'd11070, 32'd2387, -32'd14947, 32'd15368},
{32'd1998, 32'd560, 32'd7148, -32'd5111},
{-32'd3983, 32'd1587, 32'd7272, 32'd3541},
{-32'd7024, -32'd1629, -32'd16631, -32'd6105},
{32'd9251, 32'd4207, -32'd6055, -32'd712},
{-32'd11363, -32'd1412, -32'd7377, 32'd6328},
{-32'd3237, 32'd1601, 32'd12385, 32'd5109},
{32'd5855, -32'd7746, 32'd8739, 32'd3081},
{-32'd6275, 32'd2218, 32'd2405, 32'd7470},
{32'd8184, 32'd8115, -32'd12516, -32'd2903},
{-32'd1763, 32'd3392, -32'd6186, 32'd9342},
{-32'd463, 32'd1897, 32'd2834, 32'd13},
{32'd1367, -32'd2531, 32'd6687, -32'd647},
{32'd7659, -32'd10804, 32'd10382, -32'd2035},
{32'd3313, 32'd5229, -32'd11938, 32'd4469},
{-32'd2455, -32'd4149, 32'd6868, 32'd1940},
{32'd7454, -32'd770, 32'd4465, -32'd3332},
{32'd9370, 32'd3329, -32'd6634, 32'd7999},
{32'd8277, 32'd9218, -32'd4820, -32'd4243},
{-32'd1540, -32'd7954, -32'd8682, -32'd11004},
{-32'd12113, -32'd7365, 32'd3946, 32'd5987},
{32'd10572, 32'd1867, 32'd2636, 32'd8049},
{32'd3237, 32'd10242, -32'd1547, -32'd14071},
{32'd4608, 32'd10407, -32'd6147, 32'd6761},
{32'd203, 32'd1181, -32'd4015, -32'd3356},
{-32'd12770, -32'd18398, -32'd16923, -32'd2354},
{32'd2151, 32'd8072, 32'd3163, 32'd4484},
{-32'd6133, -32'd5034, -32'd6605, -32'd3722},
{-32'd4353, -32'd6022, -32'd756, 32'd3443},
{32'd5727, 32'd2289, -32'd1821, -32'd3277},
{32'd860, 32'd2787, -32'd1529, 32'd8212},
{32'd6791, 32'd5447, 32'd6144, -32'd4662},
{-32'd5146, 32'd481, 32'd4111, -32'd3034},
{32'd6175, 32'd12785, -32'd1971, -32'd14019},
{32'd6339, -32'd800, -32'd3671, -32'd1558},
{32'd2672, -32'd5311, 32'd2838, 32'd1520},
{32'd349, -32'd5219, -32'd2802, 32'd42},
{-32'd1388, 32'd5880, 32'd2828, 32'd4306},
{-32'd14131, 32'd4735, 32'd1569, -32'd1487},
{32'd1826, -32'd4876, -32'd968, -32'd6719},
{-32'd10864, 32'd9702, 32'd7095, -32'd1586},
{-32'd7511, 32'd3133, -32'd7387, 32'd4009},
{32'd438, -32'd1853, -32'd9098, 32'd3159},
{32'd1987, -32'd15327, -32'd14980, -32'd207},
{32'd3860, 32'd164, 32'd7337, -32'd9037},
{-32'd3301, -32'd13485, 32'd7513, 32'd15218},
{-32'd4027, -32'd8083, -32'd13217, -32'd895},
{32'd4688, 32'd11042, 32'd5537, -32'd791},
{-32'd7596, -32'd5648, 32'd8614, -32'd13150},
{-32'd3392, 32'd1188, 32'd11194, 32'd9140},
{-32'd4035, 32'd4498, -32'd8214, -32'd14328},
{32'd4109, -32'd5752, 32'd3420, 32'd4963},
{-32'd1973, -32'd2598, 32'd7465, -32'd1282},
{-32'd3881, -32'd3659, 32'd3753, -32'd73},
{32'd7275, 32'd3411, 32'd1819, 32'd8861},
{-32'd8213, -32'd554, 32'd223, 32'd10910},
{32'd5027, 32'd365, -32'd9017, -32'd213},
{32'd1264, -32'd1093, -32'd848, 32'd5634},
{-32'd8276, 32'd1583, -32'd3759, 32'd9391},
{32'd3338, 32'd8193, -32'd3425, 32'd3215},
{-32'd969, -32'd6878, -32'd22629, 32'd2303},
{32'd11690, 32'd2567, -32'd13933, -32'd17077},
{-32'd1708, -32'd5153, -32'd4772, -32'd7971},
{32'd5342, -32'd2102, -32'd807, 32'd6383},
{-32'd2221, -32'd5205, 32'd10573, 32'd204},
{32'd11959, 32'd23999, 32'd10539, 32'd5984},
{32'd1809, 32'd2542, -32'd6174, 32'd4199},
{-32'd5616, -32'd9339, -32'd279, 32'd6154},
{32'd147, 32'd2854, 32'd9035, 32'd3438},
{32'd4637, -32'd5549, 32'd5080, 32'd2984},
{32'd4305, -32'd14326, 32'd1623, -32'd6341},
{32'd4378, 32'd3401, -32'd5775, -32'd5639},
{-32'd5125, -32'd4509, 32'd5012, 32'd1220},
{32'd2626, 32'd8492, 32'd5343, 32'd1318},
{32'd6084, -32'd7294, 32'd10981, 32'd4846},
{32'd1343, 32'd3117, -32'd1706, 32'd2547},
{-32'd9675, -32'd11617, 32'd557, -32'd4355},
{32'd12453, -32'd3752, 32'd12681, 32'd6782},
{32'd2130, -32'd4952, 32'd4381, 32'd1684},
{32'd13935, -32'd1434, -32'd7871, 32'd6113},
{32'd5664, 32'd9270, -32'd1489, 32'd4147},
{-32'd1820, 32'd10682, 32'd6812, -32'd2236},
{-32'd10827, 32'd2434, -32'd1588, 32'd10993},
{32'd794, -32'd2650, 32'd572, -32'd5945},
{-32'd3967, -32'd7162, 32'd14414, -32'd1913},
{32'd567, 32'd1547, -32'd11269, -32'd1725},
{32'd6061, 32'd1448, -32'd8860, -32'd9207},
{-32'd4352, 32'd13697, 32'd4801, -32'd628},
{32'd4012, 32'd1407, 32'd222, -32'd1281},
{32'd7901, 32'd5378, 32'd2089, 32'd6123},
{32'd1923, -32'd384, -32'd5964, 32'd5047},
{-32'd18733, -32'd4989, -32'd6542, 32'd5419},
{-32'd5688, 32'd1883, -32'd8805, -32'd5769},
{32'd430, 32'd11623, 32'd5130, -32'd2215},
{-32'd2363, 32'd5139, 32'd9353, -32'd895}
},
{{-32'd12848, -32'd213, -32'd368, -32'd4921},
{32'd11888, -32'd7490, 32'd6264, 32'd844},
{-32'd8342, 32'd2529, -32'd2314, 32'd1111},
{32'd9102, -32'd12174, 32'd4148, 32'd7883},
{32'd564, -32'd2016, 32'd4143, -32'd7155},
{-32'd1505, -32'd1765, 32'd10277, -32'd4274},
{32'd2711, -32'd6655, -32'd12658, 32'd13826},
{32'd6110, -32'd9084, 32'd2544, 32'd6857},
{-32'd521, -32'd2625, 32'd1453, -32'd9809},
{32'd4412, 32'd5033, 32'd1345, 32'd5830},
{32'd5656, -32'd7629, 32'd7513, -32'd2383},
{32'd4615, -32'd3981, 32'd4076, 32'd5943},
{-32'd2648, 32'd5872, 32'd6711, -32'd8588},
{32'd7840, -32'd2181, -32'd8230, 32'd11691},
{-32'd7049, -32'd3064, -32'd4788, 32'd704},
{-32'd6146, -32'd9499, -32'd7928, -32'd1718},
{-32'd18733, 32'd1606, 32'd2547, 32'd7422},
{-32'd2114, 32'd1908, -32'd7610, -32'd5078},
{-32'd6693, -32'd3293, -32'd1275, 32'd10109},
{32'd638, 32'd8757, -32'd4568, 32'd7733},
{-32'd6001, 32'd17413, 32'd7453, -32'd115},
{-32'd8165, -32'd1389, -32'd5140, -32'd5634},
{-32'd7922, 32'd754, -32'd2413, 32'd235},
{32'd7730, -32'd1889, -32'd7462, -32'd1660},
{-32'd4782, 32'd9587, 32'd1218, 32'd3992},
{32'd4372, -32'd419, 32'd5627, -32'd9998},
{-32'd3398, -32'd18118, 32'd5637, 32'd533},
{32'd11265, 32'd29099, -32'd7475, 32'd883},
{-32'd4399, -32'd4173, 32'd2820, 32'd14869},
{32'd5945, -32'd9375, -32'd5625, 32'd8665},
{-32'd19203, -32'd26191, 32'd8878, -32'd7529},
{32'd4569, -32'd3224, 32'd7972, -32'd1283},
{-32'd6614, 32'd7574, 32'd12217, 32'd1285},
{-32'd113, -32'd6080, -32'd13367, -32'd8260},
{32'd8878, -32'd2347, 32'd1362, 32'd3181},
{-32'd3656, -32'd6317, -32'd1129, -32'd2795},
{32'd7920, 32'd6952, -32'd3164, 32'd1961},
{32'd6117, -32'd6856, -32'd3357, 32'd1192},
{-32'd10845, -32'd6263, 32'd274, 32'd3593},
{32'd3054, -32'd13174, 32'd6536, 32'd1489},
{32'd1632, -32'd932, -32'd429, 32'd5321},
{32'd5822, -32'd12057, -32'd5489, -32'd4573},
{32'd693, -32'd995, 32'd1634, -32'd6051},
{32'd5820, 32'd974, 32'd10759, -32'd8251},
{-32'd13577, 32'd6487, 32'd2163, -32'd8851},
{32'd5180, -32'd17414, -32'd666, -32'd7246},
{-32'd7417, -32'd8924, 32'd5430, -32'd1172},
{-32'd13428, -32'd10637, 32'd3862, -32'd1691},
{-32'd14659, 32'd8225, -32'd1159, -32'd639},
{32'd5916, -32'd3670, -32'd7935, 32'd3647},
{32'd7800, -32'd4259, -32'd982, -32'd3629},
{32'd13959, 32'd4542, 32'd1139, -32'd16478},
{-32'd3207, 32'd5926, -32'd7591, -32'd3430},
{32'd1008, 32'd12432, 32'd1221, 32'd1522},
{-32'd1473, 32'd980, -32'd3653, -32'd12215},
{-32'd7886, -32'd780, 32'd5855, -32'd8161},
{-32'd3527, 32'd7085, -32'd4579, 32'd6585},
{32'd3434, 32'd8133, -32'd2268, 32'd3596},
{32'd13283, -32'd5015, -32'd9657, 32'd7370},
{-32'd127, -32'd4260, -32'd710, 32'd7660},
{32'd7732, -32'd20380, 32'd4530, -32'd1261},
{32'd2405, 32'd6561, -32'd11866, -32'd5308},
{-32'd2265, 32'd120, -32'd4525, -32'd7013},
{-32'd4871, -32'd4425, -32'd7558, -32'd4925},
{32'd7488, 32'd17146, -32'd4960, 32'd2959},
{32'd9937, 32'd7382, 32'd8092, -32'd8035},
{32'd887, -32'd4935, 32'd8365, 32'd2198},
{32'd4594, -32'd1381, -32'd20391, -32'd11055},
{-32'd1595, -32'd4128, 32'd14234, -32'd6180},
{32'd8178, -32'd5458, -32'd723, -32'd5681},
{-32'd2642, 32'd9792, 32'd6950, 32'd2249},
{32'd18363, 32'd10406, 32'd2298, 32'd746},
{32'd10041, 32'd7463, -32'd987, -32'd4030},
{-32'd12834, 32'd5498, 32'd5240, 32'd15095},
{-32'd9757, 32'd1190, 32'd5735, 32'd9909},
{-32'd8527, -32'd5728, -32'd2447, -32'd10323},
{32'd226, -32'd13532, -32'd2399, 32'd4516},
{-32'd4880, -32'd19706, 32'd2631, 32'd4325},
{32'd5284, -32'd6567, 32'd7721, 32'd6767},
{32'd14997, 32'd4682, -32'd9920, -32'd12296},
{32'd8543, -32'd2085, -32'd3477, -32'd4233},
{32'd3821, -32'd2568, 32'd12533, 32'd3460},
{-32'd322, -32'd14999, 32'd4764, 32'd19889},
{-32'd4590, 32'd8702, -32'd6829, -32'd1486},
{32'd11789, -32'd4392, 32'd4357, -32'd2219},
{-32'd4576, -32'd1188, 32'd9225, -32'd14304},
{-32'd12872, 32'd10392, -32'd2928, 32'd4594},
{32'd2921, -32'd2571, -32'd5223, -32'd5541},
{32'd5067, -32'd3365, -32'd12639, -32'd1587},
{-32'd12855, -32'd3521, 32'd3269, 32'd8545},
{32'd2396, 32'd3788, -32'd8347, 32'd14404},
{32'd958, -32'd2491, -32'd8039, -32'd4822},
{32'd7660, 32'd7638, -32'd2510, -32'd5004},
{32'd13, 32'd16745, -32'd6892, 32'd5565},
{-32'd1457, 32'd13795, -32'd4026, -32'd2040},
{-32'd5951, -32'd4132, 32'd6545, -32'd2806},
{-32'd11077, -32'd11855, -32'd6494, -32'd1466},
{32'd4885, -32'd4466, -32'd2358, 32'd4770},
{32'd2316, 32'd3274, 32'd3147, -32'd5180},
{-32'd5723, -32'd13680, -32'd12087, 32'd2114},
{-32'd4978, 32'd5028, 32'd3906, -32'd12493},
{-32'd7090, 32'd4595, 32'd10348, 32'd6520},
{32'd13792, -32'd2658, -32'd4355, -32'd3993},
{-32'd5037, -32'd4028, -32'd3279, 32'd32},
{32'd3894, -32'd5340, 32'd15825, -32'd9988},
{-32'd13668, -32'd9475, -32'd3874, -32'd302},
{-32'd8672, 32'd5507, 32'd13005, -32'd2452},
{-32'd9332, -32'd7213, 32'd16442, -32'd3781},
{32'd11475, -32'd9698, -32'd3120, -32'd4464},
{32'd3998, 32'd3083, -32'd3644, 32'd5302},
{32'd15483, 32'd4099, -32'd10194, -32'd2855},
{-32'd515, -32'd800, 32'd148, 32'd2793},
{-32'd7891, -32'd3590, -32'd1792, 32'd10173},
{32'd9515, 32'd20226, 32'd3016, -32'd1638},
{-32'd6267, -32'd3831, 32'd1689, -32'd3712},
{-32'd2485, 32'd4058, -32'd1883, 32'd7692},
{32'd2319, 32'd5307, -32'd8727, 32'd6846},
{32'd3988, -32'd1617, -32'd7011, -32'd5885},
{32'd15668, 32'd7306, 32'd8955, 32'd4111},
{-32'd962, 32'd14773, 32'd1428, -32'd170},
{32'd6124, 32'd6206, -32'd2586, 32'd5749},
{32'd9038, 32'd7208, -32'd683, 32'd355},
{32'd5631, -32'd1235, 32'd7838, -32'd18626},
{-32'd6656, 32'd4568, -32'd3207, 32'd5893},
{-32'd9025, -32'd4059, 32'd11653, -32'd7629},
{32'd3262, 32'd14140, -32'd7769, 32'd23025},
{32'd4602, 32'd3509, 32'd1159, -32'd1882},
{32'd5851, 32'd1119, 32'd13937, -32'd2145},
{-32'd1604, -32'd13351, -32'd51, -32'd2048},
{32'd2713, -32'd10779, 32'd7343, 32'd2916},
{32'd1530, 32'd1623, 32'd3088, -32'd3023},
{32'd4795, 32'd3359, 32'd2843, -32'd947},
{-32'd8968, 32'd7075, -32'd11367, -32'd3321},
{32'd3408, -32'd4653, 32'd6209, 32'd13545},
{32'd4662, -32'd4916, -32'd769, -32'd10998},
{-32'd3877, 32'd15106, 32'd2427, 32'd2099},
{32'd6918, 32'd434, 32'd7016, -32'd7189},
{-32'd4817, -32'd9920, -32'd7644, -32'd12484},
{32'd4118, 32'd3972, 32'd8312, 32'd6660},
{-32'd3093, -32'd7401, 32'd5859, -32'd11227},
{-32'd13224, 32'd3968, 32'd8350, 32'd1315},
{-32'd3786, -32'd9462, 32'd998, -32'd3941},
{-32'd11463, 32'd10480, -32'd5411, -32'd10833},
{32'd3113, 32'd5374, 32'd13226, 32'd1976},
{-32'd2597, 32'd11576, -32'd5299, 32'd1930},
{32'd2817, 32'd13987, -32'd5841, 32'd1403},
{32'd358, -32'd8472, -32'd2913, -32'd8278},
{32'd1208, 32'd7692, 32'd7359, -32'd9274},
{32'd5480, -32'd927, 32'd4809, 32'd8529},
{-32'd2247, -32'd9314, 32'd4331, 32'd537},
{-32'd6770, 32'd6214, -32'd9260, -32'd10010},
{32'd7709, -32'd13095, 32'd8639, 32'd10208},
{32'd2540, 32'd9768, 32'd8593, -32'd14029},
{-32'd7181, -32'd5880, 32'd7852, -32'd3052},
{-32'd5182, -32'd7960, 32'd1918, -32'd3756},
{-32'd5634, 32'd5879, 32'd2182, 32'd10902},
{32'd6712, -32'd4506, 32'd5021, -32'd3408},
{32'd5908, 32'd5002, -32'd4553, -32'd3172},
{-32'd10256, -32'd328, 32'd1824, 32'd3886},
{-32'd3641, -32'd1433, 32'd11, 32'd2668},
{-32'd3931, 32'd7281, 32'd11672, 32'd3717},
{32'd6933, -32'd1382, -32'd676, 32'd6276},
{-32'd9291, 32'd13812, 32'd6041, -32'd9374},
{32'd1452, 32'd7602, -32'd5004, 32'd6692},
{32'd7415, 32'd6104, 32'd4813, 32'd17847},
{-32'd13978, 32'd4535, 32'd10490, -32'd472},
{32'd586, 32'd17123, -32'd4954, -32'd3393},
{32'd6112, 32'd7091, 32'd7096, 32'd1208},
{-32'd8174, -32'd4825, -32'd757, -32'd3137},
{32'd489, 32'd9481, 32'd432, -32'd816},
{32'd10883, -32'd4877, -32'd11023, 32'd2360},
{-32'd1851, 32'd7763, 32'd11142, 32'd5397},
{32'd4394, -32'd12053, -32'd2140, 32'd12512},
{32'd7519, -32'd314, -32'd7309, -32'd1595},
{-32'd1363, -32'd1094, 32'd6101, 32'd2518},
{-32'd11367, -32'd3704, -32'd6194, -32'd7107},
{-32'd1833, 32'd8507, 32'd2100, 32'd7040},
{32'd403, -32'd1245, 32'd11895, 32'd938},
{32'd9580, -32'd5832, 32'd6658, 32'd14056},
{-32'd12802, 32'd8414, 32'd985, 32'd2136},
{-32'd3565, 32'd3121, 32'd6704, 32'd4739},
{-32'd9115, 32'd6416, 32'd9911, 32'd3331},
{-32'd14089, -32'd4974, 32'd3049, -32'd1086},
{-32'd8352, -32'd1396, 32'd14528, -32'd1217},
{32'd8115, 32'd13958, -32'd14832, 32'd4034},
{-32'd943, 32'd3891, 32'd672, -32'd2997},
{32'd10493, 32'd98, 32'd6935, 32'd4538},
{-32'd3343, -32'd14798, 32'd12817, 32'd12714},
{32'd12569, -32'd4387, 32'd9995, 32'd3111},
{32'd2656, 32'd915, 32'd14581, 32'd605},
{-32'd1042, 32'd962, -32'd13825, -32'd9347},
{32'd2568, -32'd12513, -32'd5776, -32'd5298},
{32'd6272, -32'd2011, -32'd515, 32'd4789},
{32'd3244, -32'd3378, 32'd11583, -32'd6274},
{-32'd2604, 32'd7968, -32'd10888, 32'd8706},
{-32'd3642, 32'd2113, -32'd10513, 32'd2077},
{32'd1408, 32'd1186, 32'd3900, -32'd19596},
{32'd126, -32'd10514, 32'd1644, -32'd3775},
{-32'd10281, -32'd4840, 32'd13812, 32'd6535},
{32'd4695, 32'd4194, -32'd8922, -32'd3985},
{-32'd10194, 32'd1927, 32'd8301, -32'd1619},
{-32'd3195, -32'd3375, 32'd322, -32'd5910},
{32'd14102, -32'd13779, 32'd2073, -32'd2536},
{32'd24182, -32'd4830, 32'd13351, 32'd11067},
{-32'd2659, -32'd14504, -32'd1818, -32'd7158},
{32'd15284, 32'd10302, 32'd2881, -32'd866},
{-32'd4541, 32'd3213, -32'd5268, 32'd12671},
{32'd5372, 32'd335, 32'd850, 32'd12589},
{32'd2451, 32'd16937, -32'd7467, 32'd12130},
{-32'd9450, -32'd8704, -32'd2202, -32'd7495},
{-32'd3842, -32'd2398, -32'd4279, -32'd5494},
{-32'd14248, 32'd8872, -32'd10990, -32'd10128},
{32'd5814, 32'd3869, 32'd13332, -32'd18337},
{32'd10387, -32'd21194, 32'd1602, 32'd15579},
{-32'd11169, -32'd7046, -32'd12371, -32'd7683},
{-32'd1704, 32'd7258, -32'd6664, -32'd7720},
{32'd7334, -32'd9191, -32'd6905, 32'd3191},
{32'd407, -32'd2847, 32'd9843, -32'd3479},
{-32'd1051, -32'd2120, -32'd7450, 32'd2043},
{32'd10185, 32'd1897, 32'd1787, -32'd3798},
{-32'd9713, -32'd5249, -32'd4911, 32'd5893},
{32'd11924, -32'd7338, 32'd6312, 32'd673},
{-32'd10220, 32'd6045, 32'd2219, 32'd16156},
{-32'd6573, 32'd10522, 32'd4143, -32'd175},
{-32'd7501, -32'd5593, -32'd4912, 32'd2947},
{-32'd11794, 32'd15445, 32'd1367, 32'd8599},
{32'd4975, -32'd19893, 32'd5126, -32'd3174},
{32'd1287, 32'd2960, -32'd4818, -32'd16704},
{32'd1291, 32'd3276, 32'd7390, 32'd7546},
{-32'd319, 32'd3443, -32'd2533, 32'd6747},
{-32'd7803, 32'd3964, -32'd1776, 32'd5515},
{32'd12479, 32'd14233, -32'd2516, -32'd13846},
{-32'd4545, 32'd12925, 32'd12045, -32'd469},
{32'd12972, 32'd9699, -32'd6662, -32'd6106},
{32'd1513, 32'd12133, -32'd5913, -32'd4335},
{32'd1464, 32'd7941, 32'd7168, -32'd15041},
{32'd3249, -32'd1547, -32'd2724, 32'd7281},
{-32'd4236, 32'd4435, 32'd13185, -32'd4335},
{-32'd5493, -32'd2295, -32'd4449, 32'd2435},
{32'd8773, -32'd639, -32'd3795, -32'd2930},
{32'd2731, -32'd6262, 32'd2241, -32'd568},
{-32'd11408, 32'd3887, -32'd1047, -32'd4743},
{-32'd3930, -32'd1672, -32'd4988, -32'd1275},
{-32'd6282, -32'd2131, -32'd7003, 32'd10044},
{-32'd3867, -32'd1183, 32'd5588, 32'd6816},
{-32'd6373, -32'd4983, -32'd5962, -32'd4757},
{32'd8962, -32'd8226, 32'd3492, 32'd11628},
{-32'd1283, -32'd661, -32'd107, 32'd1480},
{-32'd14351, -32'd278, 32'd1663, 32'd14529},
{-32'd13625, -32'd2703, -32'd3637, 32'd3732},
{32'd5319, 32'd5213, 32'd4017, -32'd7523},
{-32'd2253, 32'd816, 32'd8680, 32'd397},
{32'd7073, 32'd4213, -32'd2469, 32'd1485},
{-32'd5457, -32'd1521, 32'd22473, -32'd7126},
{-32'd4895, -32'd801, 32'd6312, -32'd973},
{-32'd7115, 32'd1561, -32'd3717, 32'd4061},
{32'd1978, -32'd6547, 32'd3059, -32'd943},
{-32'd468, 32'd2169, 32'd10949, 32'd5339},
{32'd2611, -32'd713, 32'd10056, -32'd5684},
{32'd12337, -32'd5181, -32'd10734, 32'd2778},
{32'd21182, 32'd18549, 32'd3526, 32'd6096},
{-32'd2346, 32'd8980, 32'd5368, 32'd3081},
{-32'd11763, 32'd2080, 32'd2338, -32'd10439},
{32'd1137, -32'd2967, 32'd4161, 32'd13539},
{-32'd2345, -32'd3367, -32'd7328, -32'd1561},
{-32'd11895, 32'd12799, 32'd435, 32'd6198},
{32'd6475, -32'd3372, -32'd8974, 32'd1379},
{32'd6362, 32'd17461, -32'd10118, -32'd4480},
{32'd12248, -32'd1586, 32'd1153, -32'd10811},
{-32'd5458, 32'd11172, -32'd6642, 32'd3430},
{-32'd8133, -32'd5753, 32'd2149, -32'd343},
{-32'd2608, -32'd3372, 32'd3375, 32'd1974},
{-32'd7859, 32'd15815, 32'd4232, -32'd2467},
{32'd7615, -32'd239, 32'd5878, -32'd14981},
{-32'd13751, 32'd71, -32'd840, 32'd3298},
{32'd4177, -32'd11857, 32'd3468, 32'd768},
{32'd4128, 32'd5635, 32'd5337, 32'd2687},
{32'd11344, -32'd8242, -32'd8036, 32'd3690},
{-32'd2032, -32'd2999, -32'd4667, -32'd8645},
{32'd1429, -32'd9283, -32'd3901, -32'd11161},
{32'd1114, 32'd2959, 32'd22939, -32'd4758},
{32'd5289, 32'd10412, 32'd11029, -32'd2502},
{-32'd1945, 32'd709, 32'd12886, 32'd3101},
{32'd10587, 32'd3784, -32'd12851, -32'd11865},
{32'd798, 32'd3260, -32'd6668, 32'd1537},
{-32'd6919, -32'd9805, -32'd6676, 32'd14232},
{32'd7911, 32'd9815, 32'd3535, 32'd10056},
{32'd400, -32'd5048, -32'd2672, -32'd4976},
{32'd7426, -32'd4682, -32'd17490, -32'd2492},
{32'd17973, -32'd1667, -32'd4315, 32'd4797},
{32'd16055, -32'd10, -32'd1093, 32'd12173},
{32'd3361, -32'd2581, 32'd4196, 32'd6965},
{-32'd4277, 32'd7631, -32'd12933, 32'd7348},
{-32'd2338, -32'd315, -32'd3073, 32'd3432},
{-32'd14308, -32'd4303, 32'd1656, -32'd2851},
{-32'd11733, 32'd2184, -32'd6089, -32'd17963},
{-32'd9869, 32'd1585, -32'd6315, -32'd9406},
{-32'd6833, 32'd3108, 32'd4762, 32'd1554},
{32'd2251, -32'd6314, 32'd1547, 32'd16739},
{-32'd16628, 32'd3295, 32'd2887, 32'd8519}
},
{{32'd2083, -32'd3826, 32'd8333, -32'd300},
{-32'd2495, 32'd2790, -32'd8238, 32'd4172},
{-32'd3546, 32'd755, 32'd4137, 32'd6537},
{32'd3516, -32'd12, 32'd4525, 32'd4663},
{-32'd6675, -32'd11150, 32'd10239, 32'd3055},
{-32'd11554, -32'd5064, -32'd4317, 32'd3275},
{32'd9888, 32'd4763, 32'd6108, -32'd1614},
{32'd1416, -32'd3072, 32'd439, -32'd7077},
{32'd14089, 32'd4618, -32'd2023, -32'd1328},
{32'd8836, 32'd6551, 32'd13354, 32'd524},
{-32'd10345, 32'd12211, -32'd549, -32'd11308},
{32'd14271, -32'd14172, 32'd4179, -32'd3701},
{-32'd3423, 32'd5448, 32'd3155, 32'd1795},
{-32'd7385, -32'd999, -32'd3811, -32'd1198},
{-32'd636, -32'd5884, -32'd6010, 32'd3080},
{32'd7472, -32'd8759, 32'd120, 32'd6087},
{32'd4799, 32'd479, 32'd6387, 32'd1895},
{-32'd12363, -32'd5403, -32'd2023, -32'd3414},
{-32'd8607, -32'd1371, 32'd4320, 32'd2732},
{32'd3203, -32'd6506, 32'd5735, -32'd2746},
{32'd2418, 32'd10436, 32'd4942, 32'd855},
{32'd7244, -32'd4623, -32'd4346, 32'd3905},
{-32'd7649, -32'd8560, -32'd7218, -32'd2801},
{-32'd10441, 32'd2346, -32'd6622, -32'd3103},
{-32'd3038, 32'd7932, 32'd4196, -32'd1556},
{32'd5866, 32'd3986, 32'd1946, 32'd6121},
{32'd819, -32'd139, 32'd795, -32'd615},
{32'd959, 32'd2844, 32'd1668, 32'd2277},
{-32'd3305, 32'd353, 32'd268, 32'd2376},
{-32'd4061, 32'd3638, -32'd3475, 32'd2082},
{-32'd7089, 32'd903, 32'd774, 32'd4303},
{-32'd2018, -32'd5517, -32'd7841, -32'd2713},
{32'd3707, 32'd6359, 32'd9663, -32'd2001},
{-32'd5328, -32'd3866, -32'd3476, -32'd3124},
{32'd6796, 32'd5356, 32'd10442, 32'd4382},
{32'd1500, 32'd449, -32'd586, -32'd3129},
{-32'd5372, 32'd84, 32'd648, -32'd3378},
{-32'd12272, -32'd5991, -32'd726, -32'd4247},
{-32'd6126, 32'd2031, -32'd2762, -32'd1650},
{-32'd5484, 32'd3239, -32'd1899, -32'd1027},
{-32'd370, -32'd8456, 32'd3957, 32'd3441},
{32'd11058, 32'd16872, 32'd7334, -32'd1384},
{32'd1963, 32'd12931, 32'd1757, 32'd3200},
{-32'd43, -32'd3617, 32'd238, -32'd334},
{32'd305, -32'd2440, -32'd6263, -32'd7969},
{-32'd305, 32'd1809, -32'd1727, -32'd1956},
{-32'd4500, -32'd826, 32'd1058, 32'd4445},
{-32'd6329, -32'd5659, -32'd4677, 32'd1928},
{32'd1372, -32'd3129, 32'd3200, 32'd4597},
{-32'd6178, -32'd10797, 32'd3876, 32'd5331},
{32'd1509, 32'd3975, 32'd2234, -32'd128},
{32'd5741, -32'd7030, -32'd385, 32'd783},
{32'd11797, 32'd2511, 32'd6061, -32'd7341},
{-32'd4901, 32'd479, -32'd6592, -32'd2451},
{32'd5124, -32'd2342, -32'd1112, 32'd675},
{-32'd14157, -32'd5113, -32'd6601, 32'd1034},
{-32'd1607, -32'd3581, 32'd7953, 32'd373},
{-32'd12412, 32'd2275, -32'd5021, 32'd560},
{-32'd3193, -32'd2975, -32'd5643, -32'd4254},
{-32'd2263, -32'd2155, 32'd2435, 32'd3314},
{-32'd3906, -32'd222, 32'd3656, 32'd8872},
{-32'd9228, 32'd3020, -32'd3907, -32'd8774},
{-32'd5209, -32'd4424, -32'd9398, 32'd358},
{32'd8304, 32'd937, 32'd4112, -32'd380},
{-32'd11101, 32'd11127, 32'd5314, 32'd3534},
{32'd4878, 32'd13666, 32'd11156, -32'd631},
{-32'd8908, -32'd4238, 32'd1614, -32'd1047},
{-32'd368, -32'd6728, 32'd2577, 32'd6621},
{-32'd918, 32'd161, -32'd3729, -32'd5640},
{-32'd1493, -32'd853, 32'd1147, 32'd11051},
{-32'd387, -32'd1396, -32'd2671, 32'd2855},
{-32'd5043, 32'd4539, -32'd4732, -32'd5},
{-32'd2874, 32'd2914, -32'd11045, -32'd2985},
{32'd9289, 32'd5279, 32'd1769, -32'd6326},
{-32'd1167, -32'd3950, 32'd10555, -32'd4151},
{32'd4652, 32'd1606, -32'd1073, 32'd1760},
{-32'd4536, -32'd4843, -32'd10820, 32'd6607},
{-32'd6693, 32'd2711, -32'd5354, 32'd259},
{32'd5281, 32'd11817, 32'd4694, 32'd353},
{32'd11452, 32'd5904, 32'd849, -32'd1197},
{32'd1962, 32'd1986, 32'd8337, -32'd4433},
{32'd2015, 32'd14462, 32'd5348, -32'd1594},
{-32'd6391, -32'd711, 32'd4574, -32'd2291},
{32'd2696, -32'd12345, -32'd4546, 32'd429},
{32'd3739, -32'd6212, -32'd5946, -32'd1107},
{-32'd2806, 32'd4315, 32'd2933, -32'd103},
{-32'd4231, -32'd12573, -32'd5759, -32'd8489},
{-32'd7273, -32'd10958, 32'd911, -32'd2639},
{32'd23, -32'd7290, 32'd1293, 32'd2821},
{32'd2606, -32'd7139, -32'd128, 32'd3165},
{32'd1423, -32'd1897, -32'd3027, -32'd629},
{-32'd1784, 32'd1700, -32'd7654, -32'd6376},
{-32'd1985, 32'd1901, 32'd6537, -32'd853},
{-32'd754, -32'd4150, 32'd5404, 32'd1906},
{32'd5418, 32'd3469, 32'd29, -32'd5290},
{32'd5437, 32'd275, -32'd2326, 32'd136},
{32'd2182, 32'd4895, 32'd14212, -32'd249},
{-32'd2435, -32'd2927, -32'd3035, -32'd1229},
{32'd912, 32'd7849, -32'd62, -32'd248},
{32'd5790, 32'd4943, 32'd9577, 32'd4167},
{32'd5449, -32'd2433, -32'd4891, -32'd3660},
{32'd608, 32'd4809, -32'd10809, 32'd427},
{32'd1064, -32'd12340, -32'd1170, 32'd2779},
{32'd1368, -32'd3665, -32'd1716, 32'd8503},
{-32'd2667, -32'd609, 32'd5031, -32'd8995},
{-32'd4100, 32'd2557, -32'd5067, -32'd7141},
{-32'd10289, -32'd9307, -32'd2033, 32'd3285},
{-32'd5521, -32'd3182, 32'd2512, -32'd3845},
{-32'd3197, 32'd10801, 32'd845, 32'd884},
{32'd1784, -32'd12, -32'd5090, -32'd3869},
{-32'd731, -32'd3104, 32'd2176, 32'd1528},
{32'd9364, -32'd1968, 32'd6337, -32'd4391},
{32'd5332, 32'd473, -32'd2125, 32'd1501},
{-32'd2009, -32'd1888, 32'd2811, -32'd6041},
{32'd3420, -32'd1496, 32'd1652, -32'd3244},
{32'd11740, -32'd5519, 32'd73, -32'd3091},
{32'd16104, 32'd34, 32'd6726, -32'd2261},
{32'd5086, 32'd2522, -32'd4766, 32'd10819},
{-32'd3597, 32'd8467, -32'd1718, -32'd3176},
{32'd13120, 32'd5912, 32'd5717, 32'd4139},
{32'd7006, 32'd8406, 32'd6629, -32'd3982},
{32'd9489, 32'd8225, -32'd3065, 32'd1410},
{32'd1026, -32'd563, -32'd2671, 32'd3095},
{-32'd5392, -32'd3784, -32'd1782, -32'd4569},
{-32'd3979, -32'd2867, 32'd327, -32'd9388},
{32'd5972, 32'd7178, -32'd4543, -32'd5872},
{-32'd2554, 32'd259, -32'd5669, -32'd5068},
{-32'd14611, 32'd3883, 32'd2050, -32'd3895},
{32'd3289, -32'd8372, 32'd6971, -32'd458},
{32'd9075, -32'd4060, -32'd402, -32'd4240},
{32'd8149, -32'd361, 32'd4455, -32'd4886},
{32'd669, -32'd5587, -32'd9447, -32'd2822},
{-32'd6883, 32'd4394, -32'd2637, 32'd1149},
{-32'd3208, 32'd4502, -32'd910, -32'd4308},
{32'd8830, -32'd758, 32'd4251, 32'd4132},
{32'd8633, 32'd1607, -32'd4023, -32'd4704},
{32'd1444, -32'd5809, -32'd2918, 32'd80},
{-32'd5309, 32'd1690, -32'd10192, 32'd7685},
{32'd3453, 32'd6707, 32'd2408, -32'd2568},
{-32'd4775, -32'd12360, -32'd4743, -32'd1479},
{-32'd1865, 32'd1699, 32'd9591, -32'd4784},
{32'd4644, -32'd3062, -32'd1094, -32'd4094},
{-32'd2540, 32'd5144, -32'd3686, 32'd3102},
{-32'd7490, -32'd11294, -32'd4701, -32'd4173},
{-32'd333, 32'd4506, 32'd8280, 32'd2290},
{-32'd15798, 32'd3999, 32'd5293, 32'd5355},
{-32'd763, 32'd8038, -32'd630, -32'd1300},
{-32'd11301, 32'd12918, -32'd4929, -32'd3492},
{32'd8097, 32'd834, -32'd5374, 32'd454},
{-32'd5575, -32'd15644, -32'd5837, -32'd2668},
{-32'd1235, -32'd8053, -32'd8968, -32'd2148},
{32'd6700, 32'd2015, 32'd2817, 32'd4950},
{32'd3660, 32'd4533, -32'd1331, -32'd9467},
{-32'd13264, 32'd2301, 32'd3526, 32'd5590},
{-32'd6759, -32'd8269, -32'd14748, -32'd4026},
{-32'd8364, -32'd6802, -32'd301, 32'd1689},
{32'd14698, 32'd4577, -32'd272, 32'd7256},
{-32'd9366, -32'd5273, 32'd4652, -32'd5246},
{-32'd11228, -32'd1475, -32'd2943, 32'd3520},
{32'd3242, -32'd5149, 32'd3699, -32'd2437},
{-32'd11210, -32'd2380, 32'd225, 32'd7121},
{32'd3997, -32'd2231, 32'd9393, -32'd2345},
{-32'd13703, 32'd469, -32'd3135, 32'd3036},
{32'd4946, 32'd327, 32'd8021, -32'd1113},
{32'd6786, 32'd3513, -32'd4538, 32'd361},
{-32'd7009, -32'd4771, 32'd1252, 32'd1839},
{32'd5449, 32'd5984, 32'd3054, -32'd2830},
{-32'd13586, -32'd903, -32'd3245, -32'd4726},
{-32'd4535, 32'd537, 32'd5351, 32'd4707},
{-32'd5423, -32'd8081, -32'd11806, -32'd3231},
{-32'd10774, -32'd7533, -32'd13064, -32'd5420},
{-32'd12893, -32'd9192, -32'd5507, -32'd1232},
{32'd13561, 32'd1806, 32'd8067, 32'd5476},
{-32'd2464, 32'd1234, -32'd3559, -32'd7781},
{32'd8249, -32'd1964, 32'd1124, 32'd4754},
{-32'd10812, 32'd1472, -32'd1423, -32'd1539},
{32'd13587, -32'd2771, -32'd1540, 32'd32},
{32'd2000, -32'd5388, 32'd1423, 32'd4087},
{-32'd1026, -32'd13557, 32'd2815, -32'd3794},
{32'd3670, -32'd9177, -32'd6309, -32'd969},
{32'd1065, 32'd1924, -32'd2729, -32'd5906},
{-32'd5714, 32'd3422, -32'd3153, -32'd2785},
{32'd6307, 32'd3091, -32'd1457, -32'd919},
{-32'd5870, 32'd5281, -32'd3794, -32'd3385},
{32'd1656, -32'd274, 32'd2532, -32'd4272},
{-32'd2384, -32'd3558, 32'd1939, 32'd3362},
{32'd3936, 32'd652, 32'd4346, 32'd8859},
{-32'd9649, 32'd7679, -32'd308, 32'd1131},
{-32'd2144, -32'd1288, -32'd1211, 32'd2761},
{-32'd2232, -32'd2265, -32'd3788, 32'd3109},
{-32'd3581, -32'd5896, -32'd602, 32'd1058},
{-32'd5603, 32'd2255, -32'd7812, 32'd2842},
{-32'd6687, 32'd4780, -32'd4095, 32'd6566},
{-32'd7384, 32'd5264, -32'd4541, 32'd607},
{32'd17146, 32'd258, -32'd813, -32'd69},
{-32'd13369, -32'd3198, 32'd2992, 32'd73},
{32'd7605, -32'd2120, -32'd3883, 32'd1074},
{32'd1000, 32'd2441, -32'd2193, 32'd1976},
{-32'd13493, -32'd4585, 32'd3612, -32'd3754},
{-32'd3979, -32'd6297, 32'd3221, 32'd1691},
{-32'd16592, -32'd12394, -32'd9747, -32'd2589},
{-32'd2389, -32'd2664, 32'd5795, -32'd2775},
{32'd3237, -32'd3213, 32'd6090, -32'd4565},
{-32'd8637, 32'd1184, 32'd2567, 32'd5219},
{-32'd2688, -32'd9137, -32'd7224, 32'd7373},
{-32'd6775, -32'd746, 32'd2619, 32'd3423},
{-32'd2646, -32'd242, 32'd1157, -32'd920},
{-32'd1434, -32'd2779, -32'd5006, 32'd140},
{32'd4343, -32'd4688, 32'd665, 32'd3806},
{32'd14768, -32'd3121, 32'd5382, 32'd2190},
{-32'd6859, -32'd2231, 32'd1332, 32'd9460},
{-32'd4613, -32'd9342, 32'd855, -32'd5042},
{-32'd3530, -32'd4829, 32'd1078, -32'd5046},
{-32'd1284, 32'd211, 32'd3897, -32'd5075},
{-32'd2505, 32'd925, 32'd3775, -32'd3131},
{-32'd5544, -32'd9070, -32'd5405, 32'd1511},
{-32'd1717, 32'd438, -32'd3141, -32'd920},
{32'd8543, 32'd5478, 32'd3013, 32'd5233},
{32'd156, 32'd3050, -32'd1430, 32'd2609},
{32'd12205, 32'd5723, 32'd3669, -32'd1535},
{-32'd14801, -32'd12007, -32'd4478, -32'd2248},
{32'd4591, 32'd9482, 32'd5619, 32'd778},
{32'd12081, -32'd1300, 32'd4561, -32'd4001},
{32'd1129, 32'd7241, 32'd191, 32'd737},
{32'd2634, -32'd2659, 32'd323, -32'd146},
{32'd5939, -32'd9850, 32'd2216, 32'd7761},
{32'd2036, -32'd3187, -32'd967, 32'd1264},
{-32'd4480, 32'd4222, -32'd1177, 32'd119},
{32'd437, 32'd514, 32'd3970, 32'd3566},
{32'd12361, 32'd3168, 32'd7694, 32'd7137},
{-32'd8196, 32'd3446, -32'd900, -32'd1685},
{-32'd1201, 32'd5438, 32'd826, -32'd10635},
{32'd5502, 32'd1812, -32'd157, 32'd4376},
{-32'd4747, -32'd1516, 32'd4290, 32'd1481},
{-32'd5132, -32'd9001, 32'd4526, 32'd5432},
{-32'd7000, -32'd1382, -32'd2637, -32'd718},
{-32'd10078, -32'd4930, -32'd5400, -32'd5489},
{32'd10056, -32'd717, -32'd2171, 32'd2409},
{32'd14974, 32'd3208, 32'd6056, 32'd3172},
{-32'd3091, 32'd319, -32'd4807, -32'd6601},
{-32'd1270, -32'd2373, 32'd2818, -32'd2122},
{32'd3911, -32'd6321, 32'd7420, 32'd2865},
{-32'd8422, -32'd9974, -32'd11773, 32'd6438},
{32'd489, -32'd10141, -32'd5007, -32'd1223},
{32'd4472, 32'd9517, 32'd13234, -32'd2526},
{32'd11831, 32'd216, 32'd1383, -32'd6948},
{32'd567, -32'd3467, -32'd4501, -32'd7049},
{-32'd1224, -32'd6796, -32'd2369, 32'd1334},
{-32'd703, 32'd3969, 32'd735, 32'd2089},
{-32'd11723, -32'd3090, 32'd3035, 32'd7179},
{-32'd6818, 32'd10477, -32'd1620, -32'd7645},
{-32'd9105, 32'd4419, -32'd893, 32'd921},
{32'd1284, 32'd6697, 32'd2021, -32'd2237},
{-32'd8604, 32'd2733, 32'd7912, 32'd4898},
{-32'd4243, -32'd3088, -32'd5741, -32'd4826},
{-32'd14230, -32'd6475, -32'd604, 32'd3380},
{32'd455, -32'd3396, 32'd5500, -32'd698},
{32'd17136, -32'd1436, 32'd4233, -32'd1979},
{-32'd4962, 32'd1671, -32'd5110, -32'd8933},
{-32'd4709, -32'd4165, -32'd1019, -32'd1886},
{-32'd11811, -32'd1212, -32'd5246, -32'd6116},
{-32'd2580, 32'd9302, 32'd6694, 32'd1135},
{32'd4532, -32'd5818, -32'd7547, 32'd3766},
{-32'd876, -32'd2839, -32'd124, -32'd1633},
{-32'd2314, 32'd1742, -32'd1591, 32'd3758},
{-32'd11888, 32'd6214, -32'd722, -32'd7811},
{32'd2646, -32'd3597, -32'd1962, 32'd9148},
{32'd1911, -32'd154, 32'd477, -32'd1014},
{-32'd4228, 32'd3272, -32'd6716, -32'd5912},
{-32'd19597, -32'd1435, -32'd10328, 32'd4329},
{32'd4502, 32'd1467, -32'd1295, 32'd3402},
{-32'd5284, 32'd2064, 32'd4136, -32'd1063},
{-32'd6574, -32'd3934, 32'd6581, -32'd3409},
{32'd9944, 32'd2432, -32'd6702, -32'd540},
{-32'd2598, 32'd1716, -32'd1195, -32'd7048},
{-32'd4496, -32'd4116, -32'd3386, 32'd5011},
{32'd6901, 32'd8027, 32'd13544, 32'd3841},
{32'd1140, 32'd2338, 32'd2566, 32'd3548},
{32'd5777, -32'd8601, -32'd11241, -32'd1481},
{32'd9765, -32'd3265, -32'd8646, -32'd815},
{32'd1611, 32'd5771, 32'd5713, 32'd909},
{-32'd8523, 32'd3367, 32'd44, -32'd4101},
{-32'd50, -32'd1735, -32'd6294, -32'd5316},
{32'd9649, 32'd7562, -32'd4597, 32'd4810},
{-32'd9829, 32'd11609, 32'd2511, -32'd10040},
{-32'd4269, -32'd8712, -32'd5329, -32'd6299},
{32'd1202, 32'd8528, 32'd8078, -32'd4014},
{-32'd2813, -32'd5991, -32'd8287, -32'd3926},
{32'd10755, -32'd7825, -32'd5804, 32'd4560},
{32'd1030, -32'd6666, -32'd9502, -32'd4144},
{32'd8307, 32'd2459, 32'd3173, -32'd3652},
{-32'd7716, 32'd10347, -32'd2396, -32'd3903},
{32'd1539, 32'd1970, -32'd3513, 32'd4329},
{-32'd1552, -32'd5408, -32'd4628, -32'd9848},
{32'd6834, 32'd1636, -32'd11527, -32'd7424},
{32'd2181, -32'd2215, -32'd5155, -32'd2939},
{-32'd10953, -32'd1177, -32'd2130, -32'd1088},
{-32'd2281, 32'd2306, 32'd6773, -32'd3683},
{32'd15342, 32'd544, 32'd2835, 32'd5062},
{32'd6151, -32'd5196, 32'd3049, 32'd517}
},
{{-32'd5228, 32'd8892, 32'd3742, 32'd2053},
{-32'd207, -32'd17622, -32'd4447, 32'd3196},
{-32'd2267, -32'd9229, 32'd2031, 32'd12577},
{-32'd190, 32'd10586, -32'd6209, 32'd6537},
{-32'd5509, -32'd6076, -32'd8052, -32'd1160},
{32'd7083, 32'd9425, -32'd1130, 32'd10274},
{-32'd6672, 32'd9041, 32'd2577, -32'd5541},
{-32'd9648, 32'd5667, 32'd7142, 32'd2116},
{-32'd3603, 32'd4592, 32'd8484, 32'd1547},
{32'd5896, 32'd7971, 32'd6450, 32'd3373},
{-32'd2495, -32'd4777, -32'd4078, 32'd2861},
{32'd9723, -32'd965, -32'd13062, -32'd630},
{-32'd2716, 32'd2247, -32'd10030, 32'd4470},
{32'd3852, -32'd2070, -32'd1862, 32'd8463},
{-32'd10522, -32'd4864, -32'd12131, 32'd570},
{-32'd9032, -32'd3615, -32'd573, -32'd9020},
{-32'd7949, 32'd2731, -32'd5823, 32'd2143},
{32'd12296, 32'd14583, 32'd4772, -32'd4772},
{32'd5660, 32'd895, -32'd3718, -32'd6309},
{32'd1845, 32'd10042, 32'd2035, -32'd1901},
{-32'd991, -32'd13408, -32'd3267, 32'd7025},
{-32'd2797, -32'd3576, 32'd5805, 32'd6055},
{-32'd7810, -32'd6533, 32'd3244, 32'd2754},
{32'd14654, -32'd3929, -32'd3501, -32'd3289},
{-32'd4465, 32'd11453, -32'd9715, 32'd2152},
{-32'd1439, -32'd556, 32'd2290, 32'd5855},
{-32'd11409, 32'd9102, 32'd2958, -32'd1299},
{32'd22040, 32'd8538, -32'd5215, -32'd7477},
{-32'd1991, 32'd5097, 32'd3037, 32'd6926},
{-32'd3693, 32'd2638, -32'd1272, -32'd2729},
{-32'd4481, 32'd1457, -32'd7355, -32'd3555},
{32'd1368, -32'd10306, -32'd5745, -32'd1661},
{32'd3453, -32'd3358, -32'd6386, -32'd4523},
{-32'd4543, -32'd12268, -32'd6266, -32'd5653},
{32'd4877, 32'd16055, 32'd7645, 32'd826},
{-32'd9127, -32'd3949, 32'd370, 32'd4865},
{-32'd826, 32'd5182, -32'd1642, -32'd2688},
{-32'd419, -32'd1311, -32'd5506, 32'd1233},
{-32'd653, 32'd8448, 32'd860, 32'd7738},
{32'd10101, 32'd7712, 32'd1384, 32'd3094},
{-32'd10006, -32'd7468, 32'd6794, -32'd420},
{32'd11436, 32'd11207, 32'd8329, -32'd10501},
{32'd2999, 32'd6489, -32'd6928, 32'd2820},
{32'd1275, -32'd8542, -32'd11704, -32'd3802},
{-32'd8124, -32'd2694, 32'd765, -32'd1680},
{32'd573, -32'd7504, -32'd2477, 32'd2497},
{-32'd5269, -32'd5660, 32'd1996, -32'd2075},
{32'd10005, 32'd1053, -32'd11286, 32'd5283},
{-32'd10366, 32'd10674, -32'd5051, 32'd1336},
{-32'd13402, -32'd3452, -32'd2541, -32'd593},
{32'd1119, -32'd2619, -32'd12287, 32'd5431},
{32'd5426, -32'd565, 32'd4490, -32'd7106},
{32'd8494, -32'd811, -32'd3229, 32'd1167},
{-32'd5316, -32'd4166, -32'd877, 32'd2899},
{32'd6826, 32'd10860, 32'd5357, -32'd4906},
{-32'd271, 32'd1392, 32'd1945, 32'd6364},
{32'd4709, 32'd20463, 32'd6985, 32'd7021},
{-32'd8336, -32'd6615, -32'd4871, -32'd5355},
{-32'd8737, 32'd7195, 32'd880, 32'd3304},
{-32'd4051, 32'd6012, -32'd3876, 32'd7227},
{-32'd15916, -32'd7015, -32'd6083, 32'd5709},
{32'd4329, -32'd2865, -32'd1037, -32'd5640},
{-32'd7691, -32'd4713, 32'd2306, 32'd1626},
{-32'd13053, 32'd1160, 32'd5186, 32'd14676},
{32'd3933, 32'd203, -32'd9181, 32'd1649},
{32'd11581, 32'd14128, -32'd3021, 32'd1413},
{-32'd820, 32'd4018, -32'd5617, 32'd2970},
{32'd16925, 32'd2700, -32'd4483, 32'd313},
{32'd1088, -32'd8723, -32'd3873, -32'd5132},
{32'd4636, 32'd11224, 32'd12619, -32'd2965},
{32'd2514, 32'd5873, 32'd6660, -32'd6243},
{32'd5115, -32'd5073, 32'd7805, -32'd9543},
{-32'd9372, -32'd16902, -32'd587, -32'd9316},
{32'd9758, 32'd3931, -32'd1124, 32'd6805},
{32'd4148, 32'd9410, 32'd7864, 32'd6149},
{32'd14023, 32'd10639, -32'd2001, -32'd5054},
{-32'd8125, -32'd4422, -32'd11566, 32'd1375},
{-32'd425, 32'd5639, -32'd6378, 32'd11582},
{-32'd6887, 32'd6187, 32'd5363, -32'd2961},
{32'd385, 32'd5748, 32'd8230, 32'd2301},
{-32'd15495, 32'd10901, -32'd6990, -32'd3299},
{32'd4135, 32'd5425, 32'd896, 32'd1817},
{-32'd21438, 32'd3247, -32'd6948, 32'd3157},
{-32'd4026, 32'd8982, -32'd12029, 32'd3160},
{-32'd4354, -32'd13774, -32'd13309, 32'd2571},
{-32'd5143, -32'd7180, 32'd463, -32'd4452},
{32'd7897, 32'd4436, 32'd2, -32'd5107},
{-32'd7968, -32'd9733, 32'd3944, -32'd245},
{32'd1835, 32'd4491, -32'd4352, 32'd1929},
{-32'd2108, -32'd1224, -32'd2118, 32'd6488},
{32'd2366, 32'd2056, 32'd287, -32'd4394},
{-32'd6252, -32'd12885, -32'd10405, 32'd3580},
{32'd5920, 32'd8059, -32'd5604, 32'd1156},
{32'd19390, -32'd7320, 32'd11388, 32'd7169},
{32'd3333, -32'd3310, 32'd7584, -32'd7139},
{-32'd8685, -32'd4890, 32'd8812, -32'd2241},
{32'd371, 32'd15012, -32'd76, -32'd3118},
{32'd5197, 32'd6619, 32'd5486, 32'd32},
{32'd4667, 32'd7648, 32'd5606, 32'd4840},
{-32'd8277, 32'd7734, 32'd4645, -32'd6400},
{-32'd8044, -32'd6130, 32'd11402, -32'd3552},
{-32'd4240, 32'd1207, -32'd869, -32'd5883},
{32'd7213, -32'd12478, 32'd915, -32'd207},
{-32'd3389, 32'd1604, -32'd3842, 32'd4144},
{32'd1208, -32'd4529, -32'd1781, -32'd7369},
{-32'd107, 32'd5922, 32'd6681, 32'd4118},
{32'd5964, -32'd1481, 32'd4725, 32'd3523},
{-32'd5101, -32'd8589, -32'd6637, 32'd10530},
{32'd5043, -32'd1498, -32'd5982, -32'd486},
{-32'd2949, -32'd11121, 32'd8983, 32'd1785},
{-32'd12704, -32'd2582, -32'd1892, 32'd1961},
{-32'd6056, 32'd6661, 32'd9284, -32'd744},
{32'd2494, 32'd4634, -32'd5911, 32'd3232},
{32'd4959, 32'd1505, -32'd10160, -32'd4478},
{-32'd4841, -32'd13344, 32'd2174, 32'd3836},
{-32'd8004, -32'd718, -32'd6867, 32'd992},
{-32'd14069, 32'd9479, 32'd1892, 32'd2882},
{-32'd12272, 32'd3031, 32'd9452, -32'd2284},
{-32'd4385, -32'd8378, 32'd8706, -32'd5759},
{32'd14854, 32'd5650, 32'd2157, 32'd2868},
{32'd5585, -32'd9409, 32'd7280, 32'd5556},
{32'd1036, -32'd10006, 32'd3658, 32'd4649},
{32'd9842, -32'd3603, 32'd1271, -32'd3393},
{32'd7740, 32'd11277, 32'd6791, 32'd2103},
{32'd5676, 32'd3073, -32'd10401, 32'd4299},
{32'd10615, 32'd8687, 32'd8334, 32'd5287},
{-32'd6903, 32'd1784, -32'd2515, -32'd4588},
{-32'd8445, -32'd5751, 32'd5198, -32'd717},
{-32'd2167, -32'd3850, -32'd4930, 32'd811},
{-32'd2726, 32'd1765, -32'd5195, -32'd5702},
{32'd4564, -32'd2526, 32'd2261, 32'd2710},
{-32'd89, -32'd4047, -32'd8539, -32'd4329},
{-32'd6429, -32'd1504, -32'd1086, -32'd2656},
{32'd3779, 32'd17968, 32'd5417, 32'd1753},
{32'd16063, 32'd4048, 32'd2319, -32'd7468},
{-32'd3234, 32'd3189, -32'd2693, -32'd5318},
{32'd8625, 32'd7111, -32'd1301, -32'd375},
{-32'd7709, -32'd4458, -32'd1608, -32'd2252},
{32'd13669, -32'd5753, -32'd7706, 32'd2319},
{-32'd14158, 32'd1785, -32'd1753, 32'd921},
{32'd2826, 32'd9134, 32'd1924, 32'd3061},
{-32'd2324, -32'd1345, 32'd7062, -32'd1024},
{32'd14295, -32'd11457, -32'd586, -32'd2915},
{-32'd4552, -32'd9810, -32'd10355, 32'd12202},
{32'd666, 32'd1841, -32'd3001, -32'd3415},
{-32'd898, 32'd2541, -32'd6356, 32'd2489},
{-32'd561, -32'd8680, 32'd95, -32'd2501},
{-32'd14145, 32'd9331, 32'd4064, -32'd156},
{-32'd5192, 32'd1886, 32'd687, 32'd6887},
{32'd6568, -32'd9439, -32'd7375, -32'd6166},
{32'd8475, -32'd13177, -32'd9534, -32'd5502},
{32'd2167, 32'd994, -32'd2324, -32'd6702},
{-32'd4711, -32'd12243, -32'd2797, 32'd3074},
{-32'd10026, 32'd12183, 32'd3307, 32'd6120},
{-32'd1386, -32'd3725, -32'd1919, -32'd7404},
{-32'd3266, 32'd5736, -32'd7461, -32'd4061},
{32'd10036, 32'd11535, 32'd1340, 32'd2170},
{32'd18723, 32'd10141, -32'd172, 32'd2966},
{32'd1246, -32'd4565, -32'd9110, 32'd3793},
{-32'd12646, 32'd4123, 32'd3217, 32'd5277},
{-32'd14028, -32'd2782, -32'd9982, -32'd5686},
{32'd510, 32'd8139, 32'd9013, 32'd6712},
{-32'd6303, 32'd7883, -32'd6841, -32'd9401},
{32'd15645, 32'd10494, 32'd9465, 32'd8315},
{32'd7510, -32'd78, -32'd4329, 32'd8830},
{32'd3079, -32'd18594, -32'd7229, -32'd323},
{-32'd7584, -32'd9871, 32'd660, -32'd2157},
{32'd2548, -32'd140, -32'd9873, -32'd567},
{-32'd7033, -32'd4532, -32'd8745, -32'd599},
{-32'd864, 32'd3171, -32'd1551, 32'd182},
{32'd4265, 32'd4222, -32'd2724, 32'd9615},
{-32'd179, -32'd2518, 32'd325, 32'd1836},
{32'd4415, 32'd17377, 32'd7621, -32'd979},
{32'd3972, 32'd5011, -32'd2864, -32'd4170},
{32'd11031, -32'd950, -32'd5057, 32'd1729},
{-32'd5981, -32'd4311, -32'd9812, -32'd5584},
{-32'd4824, -32'd689, 32'd1571, 32'd4534},
{32'd6880, 32'd501, 32'd6016, -32'd3992},
{32'd6275, 32'd764, 32'd8663, 32'd2282},
{-32'd935, -32'd7219, -32'd14797, -32'd1498},
{32'd1066, -32'd6677, -32'd1453, -32'd5246},
{-32'd6841, -32'd8925, -32'd8822, -32'd3858},
{32'd2542, -32'd1767, -32'd12147, -32'd10228},
{-32'd10488, -32'd2330, -32'd6837, -32'd1604},
{32'd586, -32'd6390, -32'd347, 32'd3162},
{-32'd4149, 32'd5179, 32'd4488, 32'd1546},
{-32'd4412, 32'd10971, 32'd12684, -32'd705},
{-32'd4243, -32'd4673, -32'd7853, -32'd684},
{-32'd8641, -32'd9817, 32'd1378, 32'd6689},
{-32'd5229, -32'd3268, -32'd17520, -32'd12128},
{-32'd3691, 32'd4588, 32'd2608, -32'd8620},
{-32'd8115, -32'd3558, -32'd4535, -32'd3377},
{-32'd14108, -32'd3803, -32'd4488, -32'd3785},
{32'd8730, -32'd9235, -32'd431, -32'd1863},
{32'd12332, 32'd5532, 32'd1336, 32'd2786},
{-32'd1881, 32'd7421, -32'd1086, -32'd14633},
{-32'd2566, -32'd4353, -32'd2857, -32'd7749},
{32'd9887, -32'd6276, -32'd2540, 32'd1106},
{-32'd8685, 32'd9052, -32'd6390, -32'd983},
{-32'd6907, 32'd3217, 32'd5312, -32'd15521},
{-32'd5082, -32'd10863, -32'd1347, -32'd2668},
{-32'd9654, -32'd5578, 32'd10304, 32'd982},
{-32'd4943, -32'd3031, 32'd1850, -32'd2549},
{32'd11196, 32'd10355, -32'd7506, 32'd1536},
{32'd8064, 32'd2538, -32'd6264, 32'd4717},
{32'd14270, 32'd4525, 32'd8201, 32'd3632},
{-32'd11115, 32'd8019, 32'd2913, 32'd10850},
{-32'd7411, -32'd4037, -32'd15100, -32'd4409},
{32'd4835, 32'd6014, 32'd9899, 32'd167},
{32'd5314, -32'd5, 32'd3614, -32'd10906},
{32'd1328, -32'd16268, 32'd4426, 32'd1174},
{-32'd4910, 32'd1395, -32'd10697, -32'd3626},
{32'd5428, -32'd15469, 32'd1417, 32'd3202},
{-32'd2240, -32'd7712, 32'd8942, 32'd5906},
{-32'd3623, -32'd434, -32'd562, 32'd427},
{-32'd5771, 32'd2035, -32'd5451, -32'd4042},
{-32'd1862, 32'd9293, 32'd7657, 32'd16077},
{32'd8204, -32'd6893, -32'd9461, 32'd9357},
{32'd12677, 32'd18337, 32'd4618, 32'd3949},
{32'd7735, 32'd5192, 32'd101, -32'd544},
{-32'd2704, 32'd5861, -32'd2244, -32'd6329},
{-32'd3462, -32'd5595, -32'd4846, -32'd3922},
{32'd415, 32'd2948, 32'd5779, 32'd1347},
{-32'd228, -32'd514, -32'd7177, -32'd4762},
{32'd3971, 32'd2597, -32'd447, 32'd3992},
{32'd12003, -32'd2753, 32'd6384, 32'd5573},
{-32'd925, 32'd1595, -32'd3497, -32'd8},
{-32'd10974, 32'd3329, 32'd3488, 32'd1196},
{-32'd8, -32'd2383, 32'd45, -32'd4006},
{32'd3677, 32'd1060, 32'd8036, 32'd6711},
{-32'd11713, 32'd10460, 32'd9783, -32'd2904},
{-32'd865, 32'd1978, -32'd8418, -32'd3154},
{32'd2385, -32'd6581, 32'd8145, 32'd7815},
{-32'd3440, -32'd8568, -32'd3417, -32'd1152},
{-32'd1684, -32'd8581, -32'd2339, -32'd8039},
{-32'd3028, -32'd2550, -32'd1220, -32'd4100},
{-32'd2583, -32'd11379, -32'd8081, 32'd11192},
{32'd8356, -32'd3723, -32'd3436, 32'd7354},
{-32'd4512, 32'd17849, -32'd3666, -32'd9209},
{32'd151, 32'd2131, 32'd3124, -32'd4433},
{-32'd1168, -32'd5788, 32'd3882, -32'd174},
{32'd5142, 32'd693, -32'd9799, -32'd2753},
{-32'd6368, -32'd8753, -32'd5527, 32'd5570},
{-32'd6406, -32'd3467, 32'd192, 32'd9069},
{32'd5707, 32'd1608, 32'd1572, 32'd1692},
{-32'd4855, -32'd3184, -32'd1599, -32'd3467},
{-32'd4558, 32'd7059, -32'd309, -32'd3018},
{32'd806, 32'd10049, 32'd3377, 32'd4548},
{32'd7226, 32'd7973, 32'd4245, -32'd2443},
{-32'd7866, -32'd1102, -32'd339, 32'd9724},
{-32'd12889, 32'd10274, -32'd4522, 32'd3137},
{32'd8776, 32'd1486, 32'd4665, -32'd7854},
{32'd195, 32'd12795, -32'd2071, -32'd9160},
{-32'd10605, -32'd15522, 32'd1929, 32'd8229},
{-32'd5566, -32'd2053, 32'd1897, 32'd1197},
{-32'd10926, 32'd10367, 32'd8504, -32'd2955},
{-32'd122, -32'd6683, 32'd733, 32'd4200},
{32'd5311, 32'd9480, -32'd3700, 32'd1520},
{-32'd11465, -32'd3178, 32'd635, -32'd3137},
{32'd15726, 32'd3425, -32'd1313, 32'd4373},
{32'd7862, 32'd3203, 32'd11700, 32'd1177},
{32'd4887, -32'd6108, -32'd7857, -32'd4765},
{-32'd466, -32'd13732, -32'd3457, 32'd1987},
{32'd4613, 32'd365, -32'd4323, -32'd586},
{-32'd2299, -32'd515, -32'd3247, -32'd7279},
{32'd4772, 32'd7644, 32'd1702, -32'd2490},
{32'd5987, 32'd1240, 32'd4786, -32'd1275},
{32'd1010, 32'd802, -32'd952, -32'd11913},
{-32'd4129, -32'd4973, -32'd7537, -32'd7703},
{-32'd3416, 32'd2232, -32'd4557, 32'd11187},
{32'd6681, 32'd3488, -32'd6001, 32'd4521},
{-32'd1891, 32'd10733, 32'd197, 32'd5685},
{-32'd114, -32'd7318, 32'd2873, -32'd5074},
{-32'd6348, -32'd1195, -32'd4241, -32'd7925},
{32'd645, 32'd5993, -32'd9311, -32'd1997},
{-32'd426, 32'd5041, 32'd2300, 32'd10524},
{32'd4433, 32'd10291, -32'd495, 32'd3371},
{32'd7768, 32'd4610, -32'd629, -32'd8727},
{32'd90, -32'd3723, -32'd10898, 32'd2389},
{32'd6077, -32'd11252, 32'd6179, -32'd11168},
{32'd3490, -32'd8156, 32'd3645, -32'd1965},
{-32'd708, 32'd5887, 32'd7204, 32'd3621},
{32'd3808, 32'd9853, 32'd4742, 32'd11271},
{32'd4188, 32'd1944, 32'd7730, 32'd2692},
{-32'd9944, -32'd2991, -32'd3879, -32'd2235},
{-32'd5421, -32'd4676, -32'd1337, -32'd8140},
{32'd3131, 32'd12530, 32'd1924, 32'd1700},
{-32'd2306, -32'd11223, -32'd1450, -32'd2103},
{32'd13380, -32'd10107, -32'd1885, -32'd2153},
{-32'd2478, -32'd6257, -32'd1466, -32'd3431},
{-32'd1345, -32'd5660, 32'd6187, 32'd1690},
{32'd2565, 32'd5990, 32'd70, 32'd3831},
{-32'd9372, 32'd2719, 32'd2689, 32'd3562},
{32'd2431, 32'd1954, -32'd3907, -32'd2093},
{-32'd1620, -32'd11182, -32'd15907, -32'd2058},
{32'd3498, -32'd1910, -32'd3134, -32'd9780},
{-32'd9483, -32'd2422, 32'd967, -32'd3688},
{32'd1665, 32'd12941, 32'd7475, -32'd2910},
{32'd3964, 32'd13657, 32'd12769, 32'd4219},
{-32'd14193, -32'd10730, 32'd1474, -32'd643}
},
{{-32'd653, -32'd13, -32'd7491, -32'd6526},
{-32'd11554, -32'd4368, 32'd1477, -32'd6277},
{-32'd2264, 32'd7850, 32'd4551, 32'd3788},
{32'd804, 32'd1902, 32'd10278, -32'd1004},
{32'd24465, 32'd1423, 32'd772, 32'd5537},
{32'd4560, 32'd9786, 32'd4565, -32'd6309},
{32'd2435, -32'd741, 32'd770, -32'd2364},
{-32'd3538, 32'd3999, 32'd767, -32'd8979},
{-32'd6171, -32'd3239, -32'd8014, 32'd7881},
{32'd8340, 32'd16652, 32'd5030, 32'd8120},
{32'd12232, -32'd10579, 32'd6852, 32'd1648},
{-32'd168, 32'd126, -32'd5083, 32'd1577},
{32'd587, 32'd7762, 32'd9552, 32'd4208},
{-32'd2924, -32'd2204, -32'd4977, -32'd9699},
{-32'd8856, -32'd2849, -32'd11695, -32'd568},
{32'd6998, 32'd286, -32'd7524, -32'd169},
{-32'd1109, 32'd8094, 32'd605, 32'd1236},
{-32'd8909, 32'd6309, 32'd6263, 32'd1649},
{32'd4764, 32'd7798, 32'd2078, -32'd7375},
{-32'd6106, -32'd5882, -32'd3227, -32'd3621},
{32'd1109, 32'd4267, -32'd2208, -32'd3641},
{-32'd3982, -32'd5084, 32'd1, -32'd8343},
{-32'd5388, -32'd2315, -32'd11858, -32'd5129},
{32'd8462, -32'd2951, 32'd4086, 32'd2268},
{32'd554, 32'd1187, -32'd3383, 32'd7562},
{-32'd8608, -32'd5965, -32'd7633, -32'd1297},
{-32'd15309, -32'd7139, -32'd9153, 32'd8690},
{-32'd4213, -32'd1750, 32'd6872, 32'd3698},
{-32'd1671, 32'd3918, 32'd2706, -32'd2230},
{32'd922, -32'd9345, -32'd4474, 32'd2978},
{32'd5515, -32'd3281, 32'd6478, 32'd3503},
{-32'd2922, -32'd13137, -32'd11834, 32'd5746},
{32'd2252, 32'd15762, 32'd3789, 32'd323},
{-32'd6453, -32'd2130, 32'd5116, -32'd3906},
{32'd1434, 32'd13485, -32'd682, 32'd14420},
{-32'd4127, -32'd5137, 32'd5560, 32'd2141},
{32'd3205, 32'd3375, 32'd5825, 32'd8517},
{-32'd6961, -32'd1623, -32'd10552, -32'd6921},
{32'd278, -32'd7691, -32'd298, 32'd3785},
{32'd667, -32'd1397, -32'd17159, 32'd2537},
{-32'd2262, -32'd855, 32'd8701, 32'd6037},
{-32'd1855, -32'd3753, -32'd6343, 32'd8402},
{32'd1240, 32'd3189, 32'd10322, 32'd1917},
{32'd2880, -32'd2610, 32'd7390, 32'd752},
{32'd648, -32'd2859, 32'd1738, -32'd5570},
{-32'd1176, -32'd3510, 32'd7077, -32'd9302},
{-32'd8617, 32'd1938, 32'd9700, -32'd17368},
{-32'd45, -32'd2286, -32'd6970, -32'd1063},
{-32'd1290, -32'd4979, -32'd5048, 32'd2788},
{-32'd4916, -32'd5976, -32'd3795, -32'd7175},
{-32'd7969, -32'd3772, -32'd4880, -32'd818},
{-32'd5355, 32'd1826, -32'd6203, 32'd9477},
{32'd948, -32'd4790, -32'd10742, 32'd2758},
{32'd8686, -32'd7472, 32'd5095, 32'd1048},
{32'd2024, -32'd649, 32'd2192, 32'd7919},
{-32'd9046, 32'd3815, 32'd9161, -32'd9130},
{-32'd5768, 32'd7480, -32'd9289, 32'd265},
{32'd3971, 32'd1440, -32'd103, -32'd9881},
{32'd933, -32'd4491, 32'd1204, 32'd3040},
{-32'd3181, -32'd5119, -32'd1915, -32'd4980},
{-32'd1510, 32'd5885, 32'd5976, 32'd570},
{-32'd9908, -32'd10172, 32'd4613, 32'd3225},
{-32'd439, -32'd5426, -32'd5436, -32'd237},
{-32'd1641, 32'd3450, -32'd2337, -32'd3085},
{32'd8458, 32'd139, 32'd688, -32'd9798},
{-32'd5682, 32'd12038, 32'd4092, 32'd7283},
{32'd207, -32'd5158, -32'd3607, 32'd8095},
{-32'd14858, -32'd5901, 32'd6341, 32'd2483},
{32'd1978, -32'd6607, -32'd9399, 32'd1199},
{-32'd6881, 32'd2749, -32'd5629, 32'd2736},
{32'd248, -32'd11450, -32'd8595, 32'd5163},
{32'd1521, 32'd2756, -32'd6947, -32'd1992},
{-32'd1655, -32'd13023, -32'd6794, 32'd6961},
{32'd5513, -32'd920, 32'd7051, -32'd2888},
{-32'd8663, 32'd3937, -32'd1817, -32'd1348},
{-32'd1700, 32'd4245, 32'd6512, -32'd9876},
{32'd4209, -32'd1462, 32'd2677, -32'd11663},
{32'd10704, -32'd14254, -32'd3516, 32'd5471},
{32'd7283, 32'd50, 32'd9159, 32'd1561},
{32'd234, 32'd1923, -32'd6848, 32'd14648},
{32'd8786, 32'd5709, -32'd2404, -32'd4539},
{32'd13392, 32'd3384, 32'd1216, -32'd3682},
{32'd5507, 32'd3503, 32'd8502, -32'd3147},
{-32'd8021, -32'd2724, -32'd8916, 32'd5523},
{32'd1775, 32'd6106, -32'd5504, 32'd8193},
{32'd8523, -32'd5946, -32'd5080, -32'd5374},
{32'd562, 32'd4375, 32'd8345, -32'd202},
{32'd2583, -32'd9687, -32'd12883, -32'd4685},
{32'd9691, -32'd3315, -32'd2303, -32'd3741},
{32'd2369, 32'd9702, -32'd8659, -32'd10229},
{-32'd1360, 32'd3578, -32'd2217, -32'd13965},
{-32'd6073, -32'd9844, -32'd2270, -32'd4096},
{-32'd3231, 32'd6040, -32'd878, 32'd2478},
{32'd6071, 32'd7391, 32'd8263, 32'd13603},
{-32'd3058, 32'd7642, 32'd13273, 32'd3235},
{-32'd2299, 32'd2719, 32'd5685, 32'd10052},
{32'd3253, 32'd13697, 32'd15853, 32'd1817},
{32'd427, 32'd4913, 32'd35, 32'd1366},
{32'd38, 32'd1464, 32'd4759, 32'd11583},
{32'd9821, 32'd10501, -32'd941, -32'd1545},
{32'd1479, 32'd5127, 32'd3229, -32'd7657},
{-32'd5371, 32'd10726, -32'd6062, 32'd462},
{32'd1400, 32'd7677, 32'd9229, -32'd2030},
{-32'd3872, 32'd6096, 32'd5550, 32'd5782},
{-32'd4753, 32'd8161, -32'd5891, 32'd8128},
{32'd12424, -32'd8173, 32'd3696, 32'd3559},
{32'd5005, 32'd2760, 32'd642, -32'd1792},
{-32'd6181, -32'd1835, -32'd12409, 32'd5193},
{32'd9429, 32'd7612, 32'd9720, -32'd1168},
{32'd10396, -32'd4852, -32'd14381, -32'd295},
{-32'd36, -32'd4103, 32'd14569, -32'd3506},
{32'd5379, -32'd3110, -32'd5527, 32'd7006},
{32'd3213, 32'd2295, -32'd1574, 32'd2297},
{32'd4658, -32'd78, 32'd7217, 32'd1594},
{32'd4913, 32'd7517, 32'd792, -32'd3878},
{-32'd4179, -32'd11636, -32'd4978, -32'd204},
{-32'd5285, 32'd1274, -32'd6990, 32'd4442},
{-32'd1112, 32'd2215, 32'd11917, -32'd6607},
{32'd3467, 32'd141, -32'd3093, -32'd353},
{32'd3386, 32'd8170, -32'd4260, 32'd15120},
{-32'd5828, -32'd1275, 32'd4761, -32'd3991},
{32'd2733, -32'd4385, 32'd8673, -32'd268},
{-32'd10112, 32'd6950, -32'd2820, -32'd686},
{-32'd73, -32'd1708, 32'd7870, 32'd3711},
{32'd3843, 32'd6495, 32'd889, 32'd8126},
{-32'd9615, -32'd4033, -32'd14698, -32'd1565},
{32'd4301, -32'd826, -32'd13776, 32'd967},
{-32'd9765, -32'd5848, -32'd9374, -32'd4399},
{32'd3912, -32'd7406, -32'd1210, 32'd556},
{-32'd6148, -32'd2553, 32'd2363, 32'd4520},
{-32'd6201, -32'd4026, 32'd6881, 32'd3306},
{32'd12811, -32'd11802, -32'd2809, -32'd8708},
{32'd1637, -32'd4181, -32'd4251, 32'd5489},
{-32'd1377, -32'd4231, -32'd10302, 32'd1477},
{-32'd834, -32'd3057, 32'd2227, -32'd4080},
{32'd9704, 32'd7604, -32'd7872, -32'd4168},
{-32'd7613, 32'd6886, 32'd8228, 32'd10252},
{32'd3008, -32'd2427, 32'd8288, 32'd1321},
{32'd7236, 32'd8116, 32'd4228, 32'd9026},
{-32'd1180, -32'd10744, -32'd1991, 32'd796},
{32'd562, -32'd6882, -32'd4604, 32'd15080},
{32'd2933, -32'd486, -32'd1784, -32'd7359},
{-32'd7789, -32'd437, -32'd8315, 32'd5543},
{-32'd3471, -32'd6357, -32'd1805, -32'd3893},
{-32'd3309, 32'd5837, 32'd9462, 32'd12549},
{-32'd6576, 32'd2876, 32'd977, 32'd10047},
{32'd5923, 32'd2274, 32'd1430, -32'd4065},
{-32'd3899, -32'd10194, -32'd1392, -32'd3290},
{-32'd3530, 32'd9337, -32'd4965, 32'd6842},
{-32'd7771, 32'd7668, 32'd10093, -32'd7609},
{32'd2387, -32'd9825, 32'd4579, -32'd1421},
{-32'd2761, 32'd2439, -32'd2565, -32'd3696},
{32'd641, 32'd5039, 32'd1314, -32'd219},
{-32'd10528, 32'd6476, -32'd5031, -32'd5443},
{32'd609, -32'd12525, -32'd5832, -32'd13756},
{-32'd5790, 32'd3662, -32'd891, 32'd2612},
{32'd4114, 32'd11444, 32'd978, -32'd424},
{-32'd5329, 32'd3244, 32'd4807, 32'd4848},
{-32'd17043, 32'd9841, -32'd5367, 32'd2446},
{32'd7781, -32'd5288, 32'd4780, 32'd360},
{-32'd4943, -32'd12183, 32'd9898, -32'd928},
{-32'd7623, 32'd7299, 32'd4597, 32'd700},
{-32'd7491, -32'd4426, -32'd4649, -32'd1709},
{32'd3355, 32'd7428, -32'd3567, 32'd5582},
{32'd1645, -32'd403, -32'd5914, 32'd4497},
{-32'd16585, -32'd11061, -32'd5610, -32'd914},
{32'd893, 32'd2693, -32'd5189, 32'd2179},
{-32'd4032, -32'd8116, 32'd339, -32'd3689},
{-32'd87, -32'd3839, 32'd733, -32'd9313},
{32'd437, -32'd5604, -32'd9325, 32'd3416},
{-32'd5994, -32'd3511, 32'd852, 32'd6109},
{-32'd6935, 32'd5624, 32'd3383, 32'd2811},
{32'd1511, 32'd12743, 32'd2971, 32'd5816},
{-32'd1772, -32'd194, -32'd7372, 32'd1401},
{-32'd4696, 32'd5099, -32'd2753, 32'd4557},
{32'd14403, 32'd3490, 32'd6871, -32'd22},
{-32'd2777, 32'd6747, 32'd2586, 32'd109},
{-32'd13025, 32'd6853, 32'd1601, -32'd8417},
{-32'd5125, 32'd9759, -32'd1306, -32'd1862},
{32'd4642, -32'd5620, 32'd38, -32'd14629},
{-32'd14226, 32'd708, -32'd2743, 32'd1260},
{32'd9313, -32'd6420, -32'd6722, 32'd1400},
{-32'd1289, -32'd14403, -32'd1935, 32'd1615},
{32'd3403, 32'd2496, -32'd11141, -32'd7473},
{32'd4020, 32'd2377, 32'd514, 32'd6950},
{-32'd825, 32'd7577, 32'd1211, -32'd1472},
{-32'd2494, 32'd7084, -32'd382, 32'd3246},
{-32'd8871, 32'd2183, -32'd577, 32'd819},
{32'd5446, 32'd4456, -32'd7366, -32'd2415},
{32'd12237, 32'd805, 32'd96, -32'd7544},
{32'd8940, 32'd3161, 32'd3185, 32'd3928},
{32'd9509, -32'd6778, 32'd693, 32'd1936},
{32'd4746, -32'd1711, -32'd4707, 32'd2120},
{-32'd5584, 32'd4458, -32'd247, 32'd11305},
{32'd1668, -32'd264, 32'd1288, -32'd2096},
{-32'd8203, 32'd6172, 32'd8116, -32'd2183},
{-32'd3828, 32'd4075, 32'd917, -32'd1806},
{-32'd2948, 32'd3010, 32'd10377, 32'd13415},
{32'd6019, 32'd3776, -32'd7119, -32'd9177},
{-32'd14545, 32'd271, 32'd12163, -32'd4394},
{-32'd1660, -32'd13036, 32'd1497, -32'd16887},
{32'd6001, -32'd2380, 32'd2342, -32'd821},
{32'd11987, -32'd7512, 32'd1168, 32'd3470},
{-32'd5047, 32'd9699, 32'd6683, 32'd989},
{32'd13267, -32'd7084, -32'd6949, -32'd2307},
{32'd1354, -32'd8846, -32'd11113, 32'd3046},
{32'd10745, 32'd5756, 32'd8544, 32'd4696},
{-32'd5192, -32'd5385, -32'd8664, -32'd7530},
{-32'd5534, 32'd3733, 32'd2760, 32'd7323},
{32'd164, 32'd9992, 32'd7451, 32'd8673},
{32'd1974, -32'd6425, -32'd3672, -32'd2021},
{-32'd11449, 32'd394, -32'd1062, 32'd4581},
{-32'd538, -32'd12682, -32'd5648, 32'd7638},
{-32'd2819, 32'd3672, 32'd3276, 32'd4626},
{32'd6360, -32'd7209, -32'd4108, -32'd10590},
{32'd7145, -32'd11822, 32'd4463, 32'd3248},
{-32'd3032, -32'd7238, -32'd3475, -32'd5333},
{32'd1897, 32'd2377, -32'd3171, -32'd1019},
{-32'd8911, -32'd6574, 32'd10202, 32'd13127},
{-32'd5917, 32'd2427, 32'd1387, -32'd741},
{32'd1422, -32'd2931, 32'd5834, -32'd11921},
{32'd7689, 32'd3850, 32'd1863, 32'd1404},
{32'd15811, 32'd10513, 32'd2673, -32'd7937},
{-32'd8135, 32'd1004, -32'd5081, -32'd6172},
{32'd22061, 32'd9511, -32'd6529, 32'd3869},
{-32'd345, 32'd4118, -32'd11574, -32'd5802},
{32'd10591, -32'd4177, -32'd3918, -32'd6109},
{32'd6393, -32'd5126, -32'd4229, -32'd8615},
{32'd5962, 32'd12449, 32'd8639, 32'd8241},
{-32'd9169, 32'd7991, 32'd1286, 32'd6141},
{-32'd10755, -32'd4061, 32'd3569, -32'd323},
{-32'd6312, -32'd452, 32'd8, 32'd8593},
{32'd5025, 32'd1608, 32'd5888, 32'd81},
{32'd14056, 32'd11641, 32'd6006, 32'd2145},
{-32'd7984, 32'd5845, 32'd9695, -32'd12971},
{32'd932, -32'd1677, -32'd7658, -32'd20878},
{32'd5543, -32'd5398, 32'd2488, 32'd3589},
{-32'd1648, -32'd3208, 32'd3700, 32'd1037},
{-32'd2566, -32'd4089, 32'd507, -32'd7113},
{32'd5845, 32'd1705, -32'd763, 32'd2111},
{-32'd7557, 32'd3464, -32'd351, -32'd3649},
{-32'd1024, -32'd2363, 32'd44, -32'd530},
{-32'd346, -32'd8245, 32'd10011, -32'd2553},
{-32'd1239, -32'd3591, -32'd6752, 32'd8505},
{32'd794, 32'd12513, 32'd3357, 32'd5656},
{-32'd5241, 32'd3734, 32'd4866, 32'd2256},
{32'd10606, -32'd1371, -32'd12139, 32'd5572},
{-32'd7645, 32'd4794, -32'd1873, -32'd3004},
{32'd15162, 32'd16854, 32'd2239, 32'd3115},
{-32'd1592, -32'd1483, 32'd7609, 32'd6510},
{32'd9953, -32'd7166, 32'd3903, -32'd890},
{-32'd8042, 32'd13130, 32'd2858, 32'd11037},
{-32'd1130, 32'd4626, 32'd9775, -32'd8399},
{-32'd451, -32'd2764, 32'd996, 32'd2552},
{32'd4092, -32'd9060, -32'd5021, -32'd6307},
{-32'd9728, -32'd2916, -32'd2053, 32'd2697},
{32'd295, -32'd2641, 32'd225, -32'd1495},
{-32'd1662, 32'd2837, -32'd949, 32'd15159},
{-32'd990, 32'd673, 32'd2128, 32'd1422},
{-32'd5933, -32'd12466, -32'd3211, -32'd565},
{-32'd12237, 32'd1865, -32'd6235, -32'd5871},
{32'd13464, 32'd7795, -32'd9261, 32'd4738},
{32'd5926, -32'd7381, -32'd1402, -32'd1049},
{-32'd3062, -32'd2974, -32'd2042, 32'd2118},
{-32'd13940, -32'd2242, 32'd2799, -32'd2437},
{-32'd5378, -32'd8543, 32'd1041, -32'd7711},
{32'd13439, 32'd12461, -32'd98, -32'd4736},
{-32'd8528, -32'd9382, 32'd6635, 32'd7990},
{-32'd979, -32'd8570, -32'd4600, -32'd5301},
{32'd1904, -32'd619, -32'd3017, 32'd3366},
{-32'd1482, -32'd2524, -32'd364, -32'd2405},
{-32'd12884, 32'd614, 32'd6151, 32'd20068},
{32'd842, 32'd5135, -32'd12927, -32'd4075},
{-32'd535, -32'd8149, -32'd7253, -32'd282},
{-32'd723, -32'd3012, 32'd15100, -32'd6659},
{32'd7213, -32'd9041, -32'd4238, 32'd3083},
{32'd6103, 32'd17780, 32'd4443, 32'd12454},
{-32'd14284, 32'd6645, 32'd5293, 32'd6462},
{-32'd6619, -32'd2931, 32'd4515, -32'd4435},
{-32'd2676, 32'd6633, -32'd608, 32'd6988},
{-32'd6219, 32'd7501, 32'd2066, 32'd2096},
{32'd8293, -32'd5617, -32'd6294, -32'd4534},
{32'd8778, -32'd13639, 32'd3102, 32'd765},
{-32'd1703, -32'd5318, 32'd1511, 32'd10986},
{-32'd4018, 32'd2920, -32'd5028, 32'd6834},
{32'd1484, -32'd9470, -32'd5276, -32'd11620},
{-32'd1519, -32'd7153, -32'd378, 32'd1897},
{32'd3905, -32'd2798, 32'd3389, 32'd6612},
{32'd3461, -32'd3936, 32'd4868, 32'd5209},
{32'd2418, -32'd2616, -32'd6372, -32'd218},
{32'd10922, 32'd7252, -32'd975, 32'd1418},
{32'd9912, 32'd2700, 32'd4570, 32'd5328},
{-32'd738, 32'd3045, -32'd18865, 32'd2929},
{32'd12913, 32'd3467, 32'd5017, -32'd8320},
{-32'd5376, -32'd921, -32'd8110, -32'd3298},
{-32'd4951, -32'd208, -32'd7326, -32'd2394},
{32'd3642, 32'd7090, 32'd4837, -32'd10044},
{-32'd5023, -32'd190, 32'd8125, 32'd7666},
{-32'd724, 32'd4071, -32'd3243, 32'd11346},
{-32'd543, -32'd9542, -32'd5739, -32'd1897}
},
{{32'd9694, 32'd1375, 32'd8250, -32'd2223},
{32'd1853, -32'd8050, -32'd7189, -32'd2629},
{32'd13426, -32'd4005, 32'd7, -32'd5137},
{32'd7164, 32'd9034, 32'd1313, 32'd382},
{-32'd2357, -32'd2032, -32'd3348, 32'd10075},
{32'd11074, -32'd1718, -32'd3028, 32'd7180},
{32'd4473, -32'd1922, 32'd1766, 32'd7438},
{-32'd2384, 32'd1060, -32'd5004, 32'd1614},
{32'd4722, -32'd2226, -32'd4046, 32'd1053},
{32'd13134, 32'd2592, 32'd6968, 32'd9686},
{32'd923, -32'd13380, -32'd725, -32'd99},
{32'd3772, -32'd3863, 32'd1263, -32'd5111},
{32'd5195, -32'd2357, 32'd4453, 32'd3353},
{32'd895, 32'd5573, -32'd8606, -32'd304},
{-32'd7034, 32'd3356, -32'd3998, 32'd1267},
{-32'd719, 32'd1018, -32'd7590, -32'd1833},
{-32'd9193, -32'd2938, 32'd6743, 32'd1125},
{-32'd819, 32'd5506, -32'd3545, 32'd1051},
{32'd2500, 32'd1830, -32'd2625, 32'd3077},
{-32'd7462, -32'd251, 32'd7164, 32'd3211},
{32'd4228, -32'd7868, -32'd4196, -32'd6259},
{-32'd15258, 32'd2118, -32'd6608, -32'd2939},
{32'd2573, 32'd1939, -32'd244, -32'd1791},
{-32'd8392, 32'd2211, -32'd7761, -32'd7090},
{32'd2032, -32'd129, 32'd9480, 32'd2997},
{32'd2984, -32'd2047, 32'd5457, -32'd2451},
{32'd338, 32'd4313, 32'd5311, 32'd6847},
{32'd4051, 32'd5345, 32'd3413, 32'd1773},
{-32'd6812, 32'd1971, 32'd999, 32'd2676},
{32'd5116, -32'd1109, 32'd4082, -32'd4376},
{32'd2132, -32'd3108, -32'd3302, 32'd7177},
{-32'd8210, -32'd3002, -32'd9355, -32'd5638},
{-32'd627, 32'd1262, 32'd7760, 32'd8840},
{-32'd3909, -32'd1996, -32'd4227, -32'd81},
{32'd506, 32'd2173, 32'd9825, 32'd7509},
{-32'd7098, 32'd6843, 32'd2096, 32'd3536},
{-32'd3470, 32'd3671, -32'd2673, -32'd147},
{32'd6824, 32'd4431, 32'd5109, -32'd53},
{32'd318, -32'd3787, -32'd4776, -32'd1400},
{-32'd4643, -32'd8519, -32'd200, -32'd62},
{-32'd9299, -32'd126, -32'd11455, -32'd652},
{-32'd4763, 32'd3682, 32'd11106, 32'd7811},
{32'd2917, 32'd1462, 32'd4779, -32'd3056},
{-32'd4799, -32'd4962, -32'd12609, -32'd2620},
{-32'd12972, 32'd798, -32'd4085, 32'd3536},
{-32'd2870, -32'd4337, -32'd2465, -32'd1748},
{-32'd3272, 32'd6917, 32'd3406, -32'd2586},
{-32'd9753, 32'd9486, -32'd4825, 32'd438},
{32'd5587, 32'd4185, 32'd8526, 32'd12637},
{-32'd418, -32'd4751, -32'd3059, -32'd3572},
{-32'd4518, -32'd5249, -32'd7047, 32'd1981},
{32'd6321, 32'd2936, 32'd9710, 32'd7090},
{32'd421, -32'd3933, -32'd5558, -32'd11595},
{-32'd782, -32'd9223, 32'd1060, -32'd1729},
{32'd5082, 32'd2496, 32'd1063, 32'd5191},
{32'd3998, 32'd4356, -32'd6944, -32'd512},
{-32'd5027, 32'd3521, 32'd5723, -32'd1140},
{-32'd3040, 32'd575, -32'd5887, 32'd2103},
{32'd5138, -32'd9814, -32'd2614, -32'd723},
{32'd12278, 32'd5407, -32'd1688, -32'd953},
{-32'd6254, 32'd22, -32'd3580, 32'd5111},
{32'd2659, -32'd5889, -32'd770, -32'd3015},
{-32'd18662, -32'd10818, -32'd6171, -32'd1601},
{-32'd4203, -32'd1875, -32'd624, 32'd4183},
{32'd3919, 32'd126, -32'd2410, 32'd282},
{32'd7711, 32'd2818, 32'd6063, 32'd14969},
{-32'd6826, 32'd2976, 32'd700, -32'd12081},
{-32'd566, 32'd125, 32'd2950, 32'd399},
{-32'd7731, 32'd1754, 32'd3382, -32'd7350},
{-32'd11371, -32'd532, 32'd1926, -32'd1283},
{32'd8819, 32'd2692, -32'd4129, -32'd2922},
{32'd496, 32'd7557, 32'd4462, 32'd3102},
{-32'd1184, 32'd6705, 32'd681, -32'd3387},
{-32'd11891, -32'd309, -32'd3506, 32'd875},
{32'd481, 32'd1074, 32'd71, 32'd1482},
{32'd297, -32'd8303, 32'd7256, -32'd9043},
{-32'd1550, -32'd5714, -32'd8004, -32'd212},
{32'd3430, 32'd2475, -32'd7338, 32'd1097},
{32'd1121, 32'd4492, 32'd8970, 32'd7901},
{-32'd3577, -32'd1258, 32'd424, -32'd3431},
{32'd7664, -32'd6322, 32'd3295, 32'd1325},
{32'd820, -32'd10156, -32'd1452, 32'd5114},
{32'd1764, 32'd1176, -32'd8385, -32'd12268},
{32'd2075, -32'd2277, -32'd11841, -32'd7096},
{32'd2006, -32'd267, -32'd11704, -32'd190},
{-32'd5638, 32'd5695, -32'd5028, -32'd754},
{32'd3219, -32'd1688, 32'd458, 32'd1970},
{-32'd9184, -32'd3607, -32'd1087, -32'd1270},
{32'd2356, 32'd2135, -32'd2392, 32'd2967},
{32'd250, -32'd1885, -32'd2766, -32'd2309},
{-32'd810, 32'd4312, 32'd3266, 32'd7994},
{-32'd9037, -32'd1488, -32'd1634, -32'd6761},
{32'd13753, -32'd2834, 32'd10159, 32'd8236},
{-32'd736, -32'd3694, 32'd3766, -32'd4746},
{32'd786, -32'd2194, -32'd5060, 32'd360},
{-32'd1205, -32'd4508, -32'd2655, 32'd5802},
{32'd4665, 32'd4631, 32'd857, 32'd10723},
{-32'd563, 32'd61, 32'd1859, 32'd2637},
{-32'd8452, 32'd1721, -32'd4537, 32'd1649},
{32'd5290, 32'd489, 32'd6274, 32'd5017},
{32'd1465, -32'd7124, -32'd3673, 32'd5771},
{-32'd4947, -32'd6976, -32'd5327, -32'd4660},
{32'd8643, 32'd100, -32'd1740, 32'd2151},
{32'd5331, 32'd2576, 32'd10241, -32'd3006},
{32'd936, -32'd1337, 32'd2835, 32'd3128},
{32'd9015, 32'd570, -32'd9162, 32'd5886},
{-32'd835, -32'd3204, 32'd1656, -32'd3318},
{32'd3259, -32'd8801, -32'd3485, -32'd7029},
{32'd13037, -32'd8305, 32'd12193, 32'd7521},
{32'd6241, -32'd1797, -32'd5112, 32'd935},
{32'd4284, -32'd2377, -32'd1532, 32'd104},
{-32'd4669, -32'd8268, -32'd2469, -32'd5431},
{32'd3885, -32'd3083, 32'd4922, 32'd140},
{-32'd2909, -32'd233, -32'd3751, 32'd7604},
{32'd3577, -32'd2352, -32'd10748, -32'd1193},
{-32'd569, 32'd1028, -32'd1089, -32'd543},
{-32'd2098, 32'd6558, 32'd6171, -32'd2932},
{-32'd4852, 32'd1888, 32'd2186, -32'd2875},
{-32'd273, 32'd687, 32'd1965, 32'd406},
{32'd8707, 32'd6921, 32'd5340, 32'd8620},
{-32'd6026, -32'd2286, 32'd4847, 32'd4024},
{-32'd3595, -32'd1249, 32'd1363, -32'd6828},
{32'd2137, 32'd5899, 32'd5030, -32'd45},
{-32'd2100, -32'd6138, -32'd2605, -32'd5078},
{32'd5806, -32'd7774, 32'd4804, -32'd416},
{32'd13314, -32'd3559, -32'd95, -32'd14541},
{-32'd9832, 32'd3134, -32'd1300, 32'd1481},
{-32'd2348, -32'd1732, -32'd11987, -32'd6206},
{32'd1098, -32'd9707, 32'd2800, -32'd9278},
{-32'd3321, -32'd3443, -32'd7420, -32'd3532},
{-32'd78, 32'd5640, -32'd705, -32'd1103},
{-32'd1612, 32'd1033, -32'd2333, -32'd4016},
{-32'd9798, 32'd1046, -32'd9209, -32'd4115},
{32'd2582, 32'd11273, -32'd70, 32'd3391},
{32'd1620, -32'd2145, 32'd4105, 32'd1672},
{-32'd6687, -32'd5, 32'd1544, 32'd2298},
{32'd1698, -32'd418, -32'd11504, -32'd1829},
{32'd4155, -32'd612, -32'd3162, 32'd2002},
{-32'd362, -32'd7460, -32'd3686, -32'd1933},
{-32'd8792, -32'd222, -32'd7758, -32'd7036},
{-32'd4762, -32'd368, 32'd1834, 32'd145},
{32'd5773, -32'd8627, -32'd4480, 32'd4986},
{32'd3824, 32'd10748, 32'd4257, -32'd4271},
{32'd474, 32'd1470, -32'd3439, -32'd13004},
{32'd13078, -32'd988, 32'd3546, 32'd3747},
{32'd10906, 32'd1077, 32'd7947, 32'd10301},
{32'd11949, -32'd2397, -32'd2730, -32'd260},
{32'd258, -32'd1662, -32'd4710, -32'd6028},
{32'd3268, 32'd630, 32'd5711, 32'd193},
{-32'd3957, 32'd10697, -32'd5124, -32'd3583},
{-32'd10748, -32'd418, -32'd2651, -32'd6073},
{32'd6307, 32'd3976, 32'd3390, 32'd7078},
{-32'd7007, -32'd2575, -32'd10573, 32'd8103},
{-32'd2116, -32'd10096, -32'd1687, -32'd475},
{-32'd7488, -32'd7918, -32'd3491, -32'd7084},
{32'd1687, 32'd387, -32'd5900, -32'd8166},
{32'd5442, -32'd925, 32'd9191, 32'd6180},
{-32'd959, 32'd3789, 32'd1688, 32'd156},
{-32'd9644, 32'd3247, -32'd4135, -32'd4588},
{32'd14389, 32'd3488, 32'd4750, 32'd13733},
{32'd1793, 32'd1998, 32'd4283, -32'd7684},
{32'd2930, -32'd1946, 32'd8283, 32'd4393},
{-32'd112, -32'd5455, 32'd6035, 32'd1557},
{-32'd434, -32'd3777, 32'd1613, -32'd964},
{32'd4029, 32'd2983, -32'd4024, -32'd1056},
{-32'd5643, -32'd4690, -32'd4075, -32'd13068},
{32'd8940, -32'd8074, 32'd416, 32'd3000},
{-32'd370, 32'd1610, -32'd601, -32'd1441},
{32'd1180, 32'd816, 32'd4573, 32'd1637},
{-32'd11678, 32'd2870, -32'd6704, -32'd6625},
{-32'd1131, 32'd2544, -32'd10512, -32'd4948},
{-32'd102, -32'd2697, -32'd1387, 32'd654},
{32'd2954, 32'd2515, 32'd6638, 32'd5785},
{32'd2572, -32'd7615, -32'd2388, -32'd1176},
{-32'd2691, -32'd4156, 32'd2007, 32'd2764},
{-32'd128, -32'd11150, 32'd268, -32'd4943},
{-32'd4814, -32'd334, -32'd1246, 32'd792},
{32'd6531, 32'd5271, -32'd2401, 32'd5652},
{32'd2409, -32'd2911, 32'd20, -32'd6886},
{-32'd107, -32'd7158, -32'd6292, -32'd9867},
{32'd7205, 32'd2062, -32'd9306, 32'd1188},
{-32'd1016, 32'd3524, -32'd1861, 32'd1806},
{-32'd6145, 32'd2164, -32'd4410, -32'd3912},
{-32'd11358, 32'd4674, 32'd2444, 32'd4218},
{32'd881, -32'd3359, -32'd1020, 32'd4544},
{32'd11670, 32'd3657, 32'd6253, 32'd3086},
{-32'd1542, 32'd8083, 32'd5759, 32'd6691},
{-32'd7213, 32'd4437, 32'd2480, -32'd4035},
{-32'd596, -32'd5797, 32'd377, 32'd4016},
{32'd1527, 32'd2837, 32'd2113, -32'd3033},
{-32'd2919, 32'd1505, 32'd8324, 32'd861},
{-32'd3462, 32'd619, -32'd6526, -32'd3072},
{32'd12871, 32'd182, -32'd3391, -32'd6300},
{-32'd708, -32'd3571, -32'd427, 32'd5811},
{32'd720, 32'd7228, -32'd4807, 32'd499},
{32'd1117, 32'd6912, 32'd2074, 32'd12681},
{32'd4525, 32'd628, 32'd4340, 32'd4750},
{-32'd3419, 32'd1465, -32'd2173, -32'd278},
{-32'd3527, 32'd3150, -32'd605, -32'd571},
{-32'd544, 32'd3743, 32'd3905, -32'd2579},
{-32'd3826, -32'd4240, -32'd7749, -32'd5820},
{-32'd7500, -32'd7602, -32'd5285, -32'd3811},
{-32'd3451, -32'd11141, -32'd2808, 32'd3077},
{32'd9228, -32'd532, 32'd2368, 32'd10896},
{-32'd8195, -32'd2310, 32'd1769, -32'd5565},
{32'd2007, 32'd8599, -32'd5717, -32'd6737},
{32'd4512, 32'd2824, 32'd6979, 32'd9655},
{32'd296, -32'd921, -32'd5320, -32'd8628},
{32'd11188, 32'd11240, -32'd8450, 32'd943},
{-32'd784, 32'd915, -32'd75, 32'd6319},
{-32'd11877, -32'd1757, -32'd315, -32'd1560},
{32'd6938, -32'd1828, -32'd6551, 32'd4540},
{-32'd14249, 32'd3941, 32'd312, -32'd4255},
{32'd5392, 32'd677, 32'd9696, 32'd1730},
{32'd1192, -32'd12790, -32'd7647, 32'd881},
{-32'd8106, -32'd8676, -32'd2064, -32'd4449},
{32'd6708, 32'd5295, 32'd4166, -32'd1712},
{-32'd5629, -32'd2234, -32'd8933, -32'd3628},
{-32'd1296, 32'd5337, -32'd1915, -32'd463},
{-32'd8068, 32'd9265, 32'd5716, 32'd1859},
{32'd78, 32'd203, 32'd3310, -32'd6709},
{-32'd3062, 32'd105, 32'd10917, 32'd594},
{32'd4019, -32'd6656, 32'd3188, -32'd1425},
{-32'd6264, 32'd2730, 32'd59, 32'd4330},
{-32'd9158, -32'd3460, -32'd5024, 32'd3665},
{32'd965, 32'd3985, -32'd9435, 32'd6796},
{-32'd948, -32'd2364, 32'd3515, 32'd1046},
{-32'd6379, -32'd6405, -32'd1701, -32'd1422},
{-32'd6610, 32'd1006, 32'd14649, -32'd8357},
{-32'd10430, -32'd588, 32'd6228, 32'd6997},
{-32'd10715, 32'd4236, 32'd4805, 32'd4661},
{-32'd1349, 32'd268, -32'd1688, -32'd9098},
{32'd2640, -32'd2155, 32'd3634, 32'd3187},
{-32'd1500, -32'd3629, 32'd4238, -32'd373},
{-32'd2337, 32'd5238, -32'd2121, -32'd1933},
{-32'd3441, 32'd5094, -32'd5858, -32'd2828},
{32'd1790, 32'd7076, -32'd4931, 32'd900},
{-32'd1530, 32'd4182, 32'd2562, -32'd2465},
{32'd13144, -32'd941, -32'd235, 32'd1983},
{32'd1800, -32'd7139, -32'd2734, -32'd7150},
{32'd4022, 32'd114, 32'd4180, -32'd448},
{-32'd3739, 32'd3292, -32'd7133, -32'd4731},
{-32'd11882, 32'd499, -32'd8284, -32'd7304},
{32'd4135, -32'd82, -32'd6930, 32'd1753},
{32'd4705, 32'd2662, 32'd8049, 32'd9243},
{32'd443, -32'd229, 32'd1590, -32'd7491},
{-32'd3916, 32'd3890, 32'd2023, -32'd7301},
{32'd3155, 32'd1266, 32'd8247, -32'd12},
{-32'd548, 32'd4283, 32'd5165, -32'd54},
{-32'd5755, 32'd6978, -32'd6809, 32'd4228},
{32'd997, -32'd4791, -32'd2568, 32'd3083},
{-32'd7019, -32'd4393, 32'd4016, -32'd1651},
{32'd6282, 32'd4340, -32'd534, 32'd2055},
{32'd1782, 32'd3552, 32'd4372, 32'd9674},
{-32'd13106, -32'd6357, -32'd6389, -32'd3919},
{32'd796, 32'd1324, 32'd2068, -32'd3717},
{32'd4880, -32'd5877, -32'd1318, 32'd4706},
{32'd280, -32'd1481, 32'd4451, 32'd1244},
{-32'd4661, -32'd2223, -32'd5780, -32'd1699},
{32'd5213, -32'd3667, -32'd7303, 32'd2807},
{32'd8783, 32'd2838, 32'd2280, -32'd1934},
{32'd4958, -32'd5702, -32'd3599, -32'd6160},
{-32'd14456, 32'd2433, -32'd2156, -32'd10563},
{-32'd21, 32'd115, -32'd516, -32'd2621},
{32'd3980, 32'd8155, -32'd2988, 32'd868},
{32'd2396, -32'd457, -32'd3162, 32'd2768},
{32'd655, 32'd2114, 32'd574, 32'd4714},
{-32'd8043, -32'd4775, 32'd4073, 32'd5974},
{-32'd12866, -32'd4487, -32'd1430, -32'd13316},
{32'd1308, 32'd10276, -32'd2583, 32'd4205},
{32'd846, 32'd2133, 32'd6775, -32'd6367},
{-32'd1918, 32'd2023, 32'd4654, 32'd2605},
{-32'd11841, -32'd6200, -32'd853, 32'd1888},
{32'd1818, -32'd5797, -32'd4889, -32'd5663},
{32'd7982, 32'd1857, -32'd915, -32'd2861},
{-32'd12975, -32'd612, -32'd2083, 32'd1480},
{32'd8799, 32'd2990, 32'd9130, 32'd10880},
{-32'd324, -32'd3068, -32'd2592, -32'd9823},
{-32'd10789, 32'd2054, -32'd9925, -32'd5240},
{32'd6061, 32'd1254, -32'd2630, -32'd3374},
{32'd11937, -32'd2863, 32'd5027, 32'd6425},
{32'd2741, -32'd4136, 32'd2442, -32'd4030},
{-32'd1874, 32'd5506, 32'd1945, -32'd7937},
{32'd781, 32'd1757, -32'd7100, -32'd3817},
{32'd3430, 32'd2004, 32'd1036, 32'd4398},
{-32'd7557, -32'd5836, -32'd12108, -32'd8957},
{32'd9672, 32'd3484, 32'd10258, 32'd1376},
{32'd4849, 32'd973, -32'd4458, 32'd59},
{32'd3712, 32'd3641, 32'd757, 32'd987},
{-32'd5116, 32'd4098, 32'd1601, 32'd2706},
{-32'd2442, -32'd2704, -32'd1239, -32'd3892},
{32'd7437, 32'd960, 32'd9223, 32'd185},
{32'd6567, -32'd4451, -32'd4172, 32'd467},
{32'd249, -32'd4241, -32'd4852, 32'd2626},
{32'd773, -32'd5601, -32'd1068, -32'd4031},
{-32'd9854, 32'd4886, -32'd1800, -32'd502},
{32'd1709, -32'd5162, -32'd4258, 32'd2781},
{-32'd3078, -32'd1973, 32'd4302, 32'd6430},
{32'd2818, 32'd2885, 32'd539, -32'd5460},
{-32'd8855, 32'd5343, -32'd11005, -32'd333}
},
{{-32'd1478, 32'd2388, 32'd4090, 32'd7022},
{-32'd3234, -32'd7131, -32'd8594, 32'd6055},
{32'd5897, -32'd9774, 32'd4962, 32'd4014},
{32'd6764, -32'd2111, 32'd8312, 32'd6476},
{32'd17135, 32'd1607, 32'd4416, -32'd3939},
{-32'd5344, -32'd6915, 32'd1578, 32'd3159},
{-32'd5195, 32'd583, 32'd2223, -32'd3534},
{-32'd7403, -32'd386, -32'd8357, -32'd7548},
{32'd4, -32'd1704, 32'd6242, -32'd5068},
{32'd10217, 32'd8850, 32'd6764, 32'd8958},
{-32'd6722, -32'd10395, -32'd2259, -32'd2327},
{32'd2277, 32'd5980, -32'd4392, -32'd3348},
{32'd4200, -32'd5564, -32'd7042, -32'd502},
{32'd4691, -32'd9647, 32'd5334, -32'd122},
{32'd741, -32'd318, -32'd5692, 32'd1748},
{-32'd3308, 32'd1249, -32'd3127, -32'd471},
{-32'd741, 32'd600, 32'd1693, -32'd386},
{32'd1393, 32'd5770, 32'd997, 32'd46},
{32'd680, 32'd1083, -32'd2267, 32'd2251},
{32'd8536, 32'd4656, 32'd5578, 32'd1682},
{-32'd2441, -32'd6250, -32'd1162, -32'd10216},
{-32'd6919, -32'd14796, -32'd3074, 32'd1469},
{-32'd5766, -32'd1387, -32'd3013, 32'd7855},
{-32'd9907, -32'd10566, -32'd14634, 32'd1172},
{-32'd2774, 32'd3598, -32'd3152, 32'd7555},
{32'd2141, -32'd2188, 32'd3108, 32'd5968},
{-32'd10682, 32'd2989, 32'd8730, -32'd7113},
{-32'd257, -32'd3507, -32'd3805, 32'd7923},
{-32'd5081, 32'd3731, -32'd2365, 32'd985},
{32'd10073, 32'd7130, -32'd1134, -32'd4783},
{-32'd8667, 32'd1476, -32'd7636, -32'd10334},
{-32'd3709, -32'd15025, 32'd7217, -32'd9184},
{32'd3437, 32'd6924, 32'd8704, 32'd4},
{-32'd3552, -32'd2197, 32'd8257, -32'd8822},
{32'd11619, 32'd8553, 32'd1773, 32'd3612},
{-32'd5331, -32'd7532, 32'd2107, -32'd7012},
{-32'd579, 32'd2651, -32'd6533, -32'd10617},
{-32'd2374, 32'd4033, -32'd8166, 32'd1394},
{-32'd10385, -32'd890, 32'd6222, -32'd300},
{-32'd15189, 32'd31, -32'd6686, -32'd7996},
{-32'd5458, -32'd816, 32'd3492, 32'd8562},
{32'd870, 32'd2185, -32'd2289, -32'd1895},
{32'd13312, -32'd1845, 32'd6258, -32'd4448},
{-32'd2701, 32'd3128, -32'd11887, 32'd2323},
{32'd1022, -32'd2678, -32'd2278, -32'd1636},
{-32'd2460, -32'd109, -32'd4239, 32'd486},
{-32'd11399, -32'd11526, 32'd4250, 32'd7130},
{32'd229, -32'd2811, -32'd3676, -32'd3398},
{-32'd2634, 32'd6091, 32'd2414, 32'd2826},
{32'd1028, -32'd4494, -32'd9181, 32'd4424},
{32'd1472, -32'd6080, 32'd7390, 32'd8156},
{32'd751, 32'd7487, -32'd9767, -32'd3486},
{-32'd4095, -32'd12828, 32'd7567, 32'd1785},
{32'd7064, -32'd2839, -32'd7414, 32'd8181},
{-32'd2275, 32'd11595, 32'd2311, 32'd5508},
{-32'd15650, -32'd7755, -32'd1856, 32'd3383},
{-32'd6695, 32'd3009, -32'd648, -32'd1348},
{-32'd6021, -32'd6857, 32'd1286, 32'd5346},
{-32'd4965, -32'd6324, -32'd10908, -32'd6663},
{-32'd2966, 32'd2721, -32'd1704, -32'd1987},
{-32'd1340, -32'd1198, 32'd9637, -32'd11870},
{-32'd10546, -32'd863, 32'd1167, -32'd9539},
{-32'd15423, -32'd1800, 32'd865, 32'd3456},
{32'd4900, 32'd3126, 32'd5771, -32'd45},
{32'd11206, 32'd2928, 32'd664, 32'd5999},
{-32'd958, 32'd4778, 32'd7058, 32'd5243},
{32'd7661, 32'd4336, -32'd5886, -32'd5109},
{32'd2309, 32'd492, -32'd4827, 32'd11473},
{32'd3785, 32'd3713, -32'd2456, 32'd934},
{32'd2107, 32'd5021, -32'd4373, -32'd5076},
{32'd5315, 32'd3593, -32'd9891, 32'd9817},
{32'd5839, -32'd179, -32'd20117, 32'd1177},
{32'd5443, 32'd4470, 32'd5184, -32'd2720},
{-32'd11261, 32'd7446, 32'd5062, -32'd4479},
{-32'd8037, -32'd3633, 32'd5117, -32'd3023},
{32'd16701, -32'd13099, -32'd10066, 32'd16013},
{32'd2433, 32'd1286, -32'd3286, -32'd1642},
{32'd3706, 32'd4235, -32'd2604, -32'd3723},
{32'd4461, 32'd8979, -32'd5981, 32'd1141},
{32'd25, -32'd2022, -32'd10408, 32'd2306},
{-32'd210, -32'd1080, 32'd790, 32'd5560},
{-32'd1144, 32'd3406, 32'd4602, -32'd2984},
{-32'd13700, -32'd16352, -32'd300, -32'd1747},
{-32'd4514, -32'd4312, -32'd4105, 32'd130},
{32'd6969, -32'd567, -32'd8058, -32'd803},
{32'd8154, 32'd2794, 32'd6796, -32'd5372},
{-32'd10, 32'd435, 32'd7153, -32'd3964},
{-32'd1346, 32'd4782, 32'd201, -32'd8509},
{-32'd2475, -32'd5986, -32'd466, 32'd19823},
{-32'd11306, -32'd3242, 32'd7341, 32'd8316},
{-32'd1131, 32'd5364, -32'd12000, 32'd4295},
{-32'd5733, -32'd2520, -32'd3176, 32'd2394},
{32'd2636, 32'd4839, 32'd1644, 32'd8581},
{32'd8530, 32'd5629, 32'd5271, 32'd2540},
{-32'd8741, -32'd14985, 32'd2027, 32'd7694},
{32'd12946, 32'd1232, -32'd14360, 32'd512},
{32'd15204, 32'd8852, 32'd7018, 32'd345},
{-32'd477, -32'd3183, -32'd7359, 32'd3938},
{32'd326, -32'd966, 32'd2480, -32'd6920},
{32'd5094, 32'd4832, 32'd3061, 32'd11891},
{-32'd5747, 32'd2188, -32'd3830, -32'd1995},
{-32'd10239, -32'd6843, -32'd4475, 32'd10637},
{32'd7278, -32'd8050, -32'd756, 32'd6882},
{-32'd1620, 32'd3850, 32'd6018, 32'd4690},
{-32'd1799, 32'd9296, -32'd9316, -32'd4128},
{-32'd934, 32'd6982, 32'd457, -32'd10362},
{-32'd4914, -32'd8076, -32'd801, 32'd282},
{32'd13085, -32'd1369, -32'd72, 32'd1326},
{32'd5011, 32'd15538, 32'd13179, 32'd4182},
{-32'd12979, -32'd7724, -32'd9238, 32'd9530},
{32'd8242, -32'd8380, -32'd9059, 32'd870},
{-32'd2876, -32'd2959, 32'd426, 32'd443},
{32'd7147, 32'd7060, 32'd550, -32'd4703},
{32'd7925, 32'd12346, 32'd1668, -32'd8385},
{-32'd4873, -32'd3349, 32'd16776, 32'd9765},
{-32'd10382, 32'd1003, -32'd1422, -32'd10019},
{-32'd4640, -32'd3783, 32'd1879, 32'd8007},
{-32'd211, 32'd3436, -32'd3509, 32'd2881},
{-32'd5005, 32'd238, 32'd5119, -32'd8614},
{-32'd2846, 32'd5076, 32'd5687, 32'd4522},
{32'd4568, 32'd847, 32'd2353, 32'd3468},
{32'd2360, -32'd3116, -32'd3655, -32'd9712},
{32'd4650, 32'd418, 32'd384, 32'd4978},
{32'd5370, -32'd580, -32'd2611, 32'd4970},
{32'd5566, -32'd3439, -32'd83, 32'd778},
{-32'd8834, -32'd6295, 32'd7539, 32'd3566},
{-32'd5893, -32'd6468, -32'd155, -32'd1121},
{32'd169, -32'd9154, -32'd13467, -32'd626},
{-32'd5346, -32'd3822, -32'd4728, -32'd9532},
{32'd657, -32'd2495, -32'd7367, -32'd9547},
{32'd1560, -32'd4154, 32'd13976, -32'd4187},
{-32'd8008, -32'd11799, -32'd11428, -32'd3909},
{-32'd10447, -32'd11548, 32'd145, -32'd9003},
{-32'd4503, -32'd4322, 32'd7384, 32'd3642},
{32'd8514, 32'd2453, 32'd311, 32'd1724},
{-32'd12345, 32'd6371, -32'd9496, -32'd5527},
{-32'd2159, 32'd7355, -32'd4619, -32'd545},
{32'd3207, 32'd3259, -32'd198, 32'd1259},
{32'd7723, -32'd2058, -32'd1268, -32'd9719},
{-32'd10141, 32'd5107, -32'd7248, -32'd3620},
{32'd5923, 32'd11033, 32'd4302, -32'd6655},
{-32'd3652, 32'd4478, -32'd5819, 32'd1762},
{32'd4249, -32'd6640, 32'd2980, -32'd801},
{-32'd8837, -32'd10078, -32'd970, -32'd6286},
{32'd7636, 32'd1829, 32'd5935, 32'd1208},
{-32'd1229, 32'd9860, 32'd510, -32'd1936},
{-32'd6735, -32'd6069, -32'd4577, -32'd12188},
{-32'd7999, 32'd7142, -32'd13084, -32'd1793},
{32'd4360, -32'd1868, 32'd5027, 32'd7637},
{-32'd4286, -32'd7971, 32'd9193, -32'd4861},
{-32'd4475, -32'd2000, -32'd12573, -32'd6429},
{32'd10675, -32'd3528, 32'd1916, -32'd2234},
{-32'd7111, 32'd2449, 32'd4063, -32'd1110},
{-32'd96, -32'd9487, 32'd2615, 32'd3748},
{-32'd10980, 32'd1916, -32'd9487, -32'd7907},
{-32'd10746, -32'd7171, 32'd2833, -32'd1997},
{32'd1599, 32'd1251, 32'd4397, 32'd12003},
{32'd597, 32'd1043, -32'd2118, -32'd671},
{32'd5720, -32'd4709, 32'd4141, -32'd4614},
{-32'd9093, 32'd17010, 32'd2851, -32'd969},
{-32'd3479, -32'd11285, -32'd21, -32'd6109},
{-32'd4802, -32'd3524, 32'd898, 32'd6459},
{-32'd7986, 32'd666, -32'd2540, -32'd1555},
{32'd7978, 32'd9326, -32'd11956, -32'd8887},
{-32'd10407, 32'd7206, -32'd2288, 32'd4336},
{-32'd2652, 32'd1176, -32'd836, -32'd2135},
{32'd1443, 32'd11460, 32'd2674, 32'd6803},
{32'd3048, -32'd1257, -32'd10651, -32'd9440},
{32'd2453, -32'd10210, 32'd3764, -32'd1595},
{-32'd7312, 32'd4785, -32'd6468, -32'd9096},
{-32'd7687, -32'd4251, 32'd1357, -32'd15000},
{-32'd15609, -32'd3647, 32'd8376, -32'd9213},
{32'd8203, 32'd5843, 32'd2370, 32'd3521},
{32'd554, 32'd522, 32'd9732, -32'd4482},
{-32'd998, -32'd6938, 32'd6737, 32'd2010},
{-32'd4076, 32'd3946, -32'd12862, -32'd8352},
{32'd7419, -32'd1378, 32'd5373, 32'd236},
{-32'd392, -32'd2181, -32'd80, 32'd7379},
{32'd5334, -32'd4133, -32'd5143, 32'd2655},
{-32'd18201, -32'd4321, -32'd7661, 32'd5041},
{32'd7, -32'd424, -32'd3449, -32'd5264},
{-32'd2100, -32'd4674, -32'd1405, -32'd7440},
{32'd6250, 32'd1180, -32'd14589, -32'd5741},
{32'd698, -32'd3149, -32'd2038, 32'd3766},
{32'd374, 32'd924, -32'd5955, -32'd2078},
{32'd5048, 32'd16683, 32'd7582, 32'd6072},
{32'd3318, 32'd594, 32'd2486, 32'd337},
{32'd3544, -32'd12089, -32'd4378, -32'd6685},
{32'd6394, -32'd3315, -32'd925, 32'd1423},
{-32'd10649, -32'd2421, -32'd3772, 32'd8605},
{-32'd3898, 32'd3701, 32'd383, -32'd1718},
{32'd4882, 32'd5303, -32'd2058, -32'd5292},
{-32'd700, -32'd7361, -32'd6556, 32'd2051},
{-32'd7857, -32'd1476, 32'd16240, -32'd603},
{32'd3764, 32'd8124, -32'd1543, -32'd1135},
{-32'd4687, 32'd9524, -32'd180, -32'd5188},
{32'd2719, 32'd10688, 32'd1928, -32'd1860},
{32'd9016, 32'd1595, -32'd6683, -32'd3620},
{-32'd12594, -32'd5761, 32'd3755, 32'd4621},
{32'd1864, 32'd16535, 32'd1002, -32'd1397},
{-32'd8619, -32'd6762, -32'd7656, -32'd3338},
{-32'd11858, 32'd11009, 32'd73, -32'd5371},
{32'd5607, 32'd2804, 32'd5509, -32'd3851},
{32'd5350, 32'd5919, 32'd7846, 32'd4582},
{32'd8052, -32'd7377, 32'd3008, -32'd4754},
{32'd4772, 32'd8562, -32'd7191, -32'd5008},
{-32'd8131, 32'd7873, -32'd1562, 32'd1125},
{32'd3391, -32'd134, -32'd10253, -32'd1712},
{-32'd4438, 32'd806, -32'd1856, 32'd13605},
{32'd3608, 32'd2529, 32'd11707, 32'd1634},
{32'd4701, -32'd2758, -32'd10063, -32'd12485},
{-32'd3912, 32'd3131, 32'd3089, 32'd1580},
{32'd2511, -32'd1276, -32'd5068, -32'd2662},
{32'd6205, 32'd2553, 32'd9818, -32'd2276},
{-32'd7552, 32'd211, 32'd296, 32'd530},
{32'd6678, -32'd4439, -32'd4680, 32'd3417},
{32'd5703, 32'd4715, 32'd3795, -32'd9237},
{-32'd2208, -32'd997, 32'd3779, 32'd8121},
{32'd3451, 32'd15935, 32'd5737, -32'd12653},
{-32'd56, -32'd3259, -32'd867, 32'd6001},
{-32'd3997, 32'd3959, -32'd3318, 32'd2283},
{32'd9588, -32'd9193, 32'd1892, 32'd548},
{-32'd1974, -32'd976, 32'd5618, 32'd8589},
{32'd765, 32'd8031, -32'd14631, 32'd9181},
{-32'd9451, 32'd1933, -32'd2655, 32'd759},
{-32'd483, -32'd5207, -32'd3294, -32'd8624},
{32'd235, -32'd6829, -32'd993, 32'd14975},
{32'd4353, -32'd2485, -32'd1670, -32'd6525},
{32'd294, -32'd9527, -32'd3, 32'd3563},
{-32'd17640, -32'd5440, -32'd4428, 32'd7591},
{-32'd7385, 32'd7344, -32'd1494, -32'd2690},
{32'd1053, 32'd3438, 32'd2294, -32'd2496},
{-32'd14983, -32'd2819, -32'd7152, -32'd201},
{32'd8345, -32'd919, -32'd1248, -32'd1336},
{32'd4922, -32'd5852, -32'd4654, 32'd6644},
{-32'd599, -32'd2955, 32'd280, -32'd4619},
{32'd813, -32'd9412, 32'd843, -32'd478},
{32'd787, -32'd15137, -32'd35, -32'd3597},
{-32'd706, 32'd5186, -32'd5154, 32'd5421},
{32'd4458, -32'd4368, 32'd566, -32'd1875},
{-32'd5225, -32'd337, -32'd180, -32'd3217},
{32'd2132, -32'd1029, 32'd4777, 32'd5342},
{-32'd18017, -32'd9355, -32'd7074, -32'd9265},
{-32'd6127, 32'd2796, 32'd8116, 32'd9676},
{32'd6354, 32'd3096, 32'd2040, 32'd5979},
{32'd13087, 32'd2959, 32'd4663, -32'd9820},
{-32'd10164, -32'd919, 32'd227, -32'd4444},
{-32'd8411, 32'd766, 32'd1663, 32'd7803},
{-32'd4751, -32'd292, -32'd6522, 32'd225},
{-32'd5685, -32'd5485, 32'd417, 32'd7736},
{-32'd7267, 32'd1403, -32'd1749, -32'd3612},
{32'd4704, 32'd1316, 32'd4972, 32'd804},
{32'd10776, 32'd4476, 32'd196, 32'd3530},
{-32'd2416, -32'd420, 32'd8967, 32'd3443},
{-32'd4738, 32'd729, -32'd8161, -32'd3236},
{-32'd8236, -32'd2117, 32'd4542, 32'd8314},
{32'd6417, 32'd2389, -32'd1607, -32'd3469},
{32'd6905, 32'd3872, 32'd678, 32'd2658},
{-32'd5850, -32'd6573, -32'd6754, -32'd10078},
{-32'd1377, 32'd2256, 32'd11284, -32'd3590},
{-32'd6005, 32'd2834, -32'd5376, 32'd3215},
{32'd7473, 32'd269, -32'd3163, -32'd4583},
{32'd3537, -32'd5187, 32'd1812, -32'd12502},
{-32'd2304, 32'd4984, -32'd6035, -32'd6943},
{32'd9284, -32'd982, -32'd10983, 32'd4632},
{-32'd9818, 32'd6038, -32'd597, 32'd18493},
{32'd1104, 32'd948, 32'd137, 32'd5898},
{-32'd1846, 32'd3782, -32'd9333, -32'd2003},
{32'd5647, -32'd13110, -32'd3294, -32'd7042},
{32'd137, -32'd3586, 32'd3246, 32'd8570},
{-32'd5748, 32'd3408, -32'd7660, -32'd890},
{32'd1151, -32'd4802, 32'd718, 32'd1866},
{-32'd9204, -32'd1505, -32'd3772, -32'd1478},
{-32'd1723, 32'd3436, -32'd1022, -32'd5833},
{-32'd3069, 32'd3340, -32'd3136, 32'd9919},
{32'd2382, -32'd3682, -32'd9985, -32'd10115},
{32'd9497, 32'd11134, 32'd6791, 32'd6488},
{-32'd527, 32'd1730, 32'd14068, 32'd7779},
{-32'd8195, 32'd2164, 32'd6772, -32'd6175},
{-32'd2605, 32'd1310, 32'd7133, -32'd5362},
{-32'd8273, 32'd6777, 32'd3390, -32'd8496},
{32'd804, 32'd8871, -32'd8325, 32'd1113},
{32'd707, 32'd3168, -32'd5381, -32'd8606},
{-32'd2671, -32'd3611, 32'd3776, 32'd5077},
{-32'd272, -32'd6436, 32'd1428, -32'd4671},
{-32'd5184, -32'd14087, 32'd3363, -32'd5486},
{-32'd2090, 32'd1951, 32'd9933, 32'd12207},
{32'd1795, -32'd3180, -32'd2162, 32'd2895},
{32'd1734, 32'd9589, 32'd8271, 32'd1930},
{-32'd7693, -32'd1931, -32'd6819, 32'd736},
{32'd4319, -32'd8246, -32'd2560, -32'd3874},
{32'd11322, 32'd1905, 32'd453, -32'd2544},
{-32'd6398, -32'd4143, 32'd821, 32'd11797},
{32'd6871, 32'd3505, -32'd6431, 32'd7101},
{-32'd8463, -32'd491, -32'd11236, 32'd1716},
{-32'd4066, 32'd4140, -32'd8799, -32'd3941},
{32'd4455, -32'd144, 32'd4355, -32'd2193},
{32'd4068, 32'd6072, 32'd8061, 32'd3357},
{-32'd798, -32'd187, 32'd15577, 32'd6687},
{-32'd6101, -32'd4023, 32'd1985, -32'd3516}
},
{{32'd10302, -32'd2932, 32'd6547, 32'd7158},
{-32'd1288, -32'd2908, -32'd574, -32'd6387},
{-32'd14087, -32'd8467, -32'd7168, -32'd1693},
{32'd13152, -32'd4475, 32'd5877, 32'd5244},
{-32'd17058, -32'd5832, -32'd6105, 32'd3572},
{-32'd5997, 32'd1450, 32'd3468, 32'd4192},
{-32'd9341, 32'd3176, 32'd2106, 32'd1193},
{32'd1717, -32'd1724, -32'd2737, -32'd1841},
{32'd5450, -32'd3002, -32'd5609, -32'd7629},
{32'd690, 32'd5110, 32'd5342, 32'd8164},
{-32'd8088, -32'd10246, -32'd3102, -32'd1257},
{32'd4572, 32'd3705, 32'd1052, 32'd6465},
{32'd13293, 32'd2111, 32'd2265, 32'd3185},
{-32'd4306, -32'd4975, -32'd116, 32'd3339},
{-32'd7863, -32'd5436, 32'd1007, -32'd4907},
{32'd1973, -32'd2308, -32'd5023, -32'd865},
{32'd22285, -32'd4946, -32'd2400, -32'd3090},
{32'd2295, -32'd8991, 32'd5943, -32'd597},
{-32'd7263, 32'd2648, -32'd3600, 32'd3712},
{-32'd7616, -32'd14556, 32'd5, 32'd5644},
{32'd465, -32'd13155, -32'd5810, -32'd520},
{-32'd2422, 32'd1660, -32'd798, -32'd2936},
{-32'd11680, -32'd12742, -32'd3225, 32'd1126},
{32'd2252, 32'd6931, -32'd15586, -32'd7352},
{-32'd543, 32'd3908, -32'd904, 32'd2710},
{32'd6021, 32'd8888, -32'd105, -32'd2391},
{32'd11464, 32'd1153, 32'd457, -32'd9386},
{-32'd1823, -32'd5372, -32'd2666, -32'd3455},
{-32'd190, 32'd5563, 32'd2414, 32'd6834},
{-32'd3105, -32'd11745, 32'd386, -32'd1109},
{-32'd2046, -32'd578, 32'd3716, -32'd1276},
{-32'd1835, 32'd10590, -32'd8225, -32'd7256},
{32'd5897, -32'd1931, 32'd12246, 32'd4152},
{32'd14987, -32'd9724, -32'd3631, -32'd4335},
{32'd4320, -32'd2542, 32'd6359, 32'd9866},
{32'd3768, 32'd8189, 32'd1348, -32'd3765},
{32'd11678, 32'd1448, 32'd1901, 32'd3372},
{-32'd1456, -32'd5146, 32'd175, 32'd4117},
{32'd2079, -32'd536, 32'd3469, 32'd1984},
{32'd6147, 32'd468, -32'd7983, 32'd637},
{-32'd4289, 32'd1399, 32'd597, -32'd4689},
{32'd401, 32'd4321, 32'd472, 32'd215},
{-32'd7722, -32'd11960, -32'd3485, 32'd1686},
{32'd271, 32'd6186, -32'd7857, -32'd3288},
{32'd8709, -32'd6211, 32'd6102, -32'd913},
{-32'd2400, -32'd680, -32'd6379, 32'd2355},
{-32'd16705, 32'd4419, -32'd1219, -32'd3753},
{32'd5722, 32'd2846, -32'd8781, -32'd1903},
{-32'd14845, -32'd1794, 32'd8174, -32'd1516},
{-32'd4855, 32'd8346, 32'd4015, -32'd46},
{32'd7591, -32'd7237, 32'd3283, 32'd4593},
{-32'd1381, 32'd5576, -32'd1499, 32'd2259},
{32'd7103, -32'd6313, 32'd1491, -32'd2779},
{32'd3379, 32'd3017, 32'd2987, -32'd1094},
{32'd1706, -32'd2218, -32'd3976, -32'd1419},
{-32'd4607, -32'd5863, -32'd3378, 32'd2618},
{-32'd11205, 32'd5500, 32'd113, -32'd90},
{-32'd1746, 32'd3795, -32'd10676, 32'd1271},
{-32'd5830, -32'd7677, 32'd2999, -32'd4587},
{-32'd6326, -32'd3806, 32'd4744, 32'd489},
{-32'd673, 32'd8245, -32'd5049, -32'd1050},
{32'd21810, -32'd4060, 32'd5472, -32'd18},
{-32'd8920, 32'd3002, -32'd5428, -32'd2609},
{-32'd4866, -32'd10686, 32'd328, 32'd271},
{-32'd8579, -32'd2073, 32'd2598, -32'd3854},
{-32'd5964, -32'd1499, 32'd3026, 32'd1991},
{32'd11456, -32'd2901, -32'd4579, 32'd1439},
{-32'd8321, -32'd11223, 32'd1214, -32'd5477},
{-32'd1642, 32'd11898, 32'd811, -32'd67},
{32'd348, 32'd4701, -32'd7204, 32'd1341},
{32'd3840, 32'd4786, -32'd8038, 32'd916},
{32'd14669, 32'd3005, -32'd6163, -32'd4862},
{-32'd2275, 32'd4388, -32'd3982, 32'd1782},
{32'd260, -32'd868, -32'd7699, -32'd4632},
{-32'd626, -32'd9854, 32'd1006, 32'd5897},
{32'd16879, 32'd909, -32'd6700, -32'd2530},
{-32'd4130, -32'd3419, -32'd6679, -32'd3204},
{32'd8283, -32'd4759, -32'd1427, 32'd2648},
{32'd4296, 32'd2312, 32'd8280, -32'd6755},
{32'd14369, -32'd427, -32'd7514, 32'd1319},
{32'd1938, 32'd4996, 32'd305, 32'd103},
{32'd11171, 32'd4611, 32'd8679, -32'd678},
{-32'd4649, 32'd6002, -32'd10718, -32'd4079},
{-32'd2980, -32'd3775, -32'd2800, -32'd1674},
{32'd3176, 32'd3255, -32'd4958, 32'd1774},
{-32'd4495, 32'd8323, -32'd5380, 32'd288},
{-32'd4494, 32'd11387, 32'd15196, 32'd5210},
{-32'd6603, 32'd1034, -32'd2744, -32'd4210},
{32'd9486, -32'd5519, 32'd3763, -32'd4588},
{32'd5856, 32'd213, -32'd8391, -32'd2042},
{-32'd4443, 32'd10356, 32'd10647, 32'd2635},
{-32'd15762, 32'd11747, -32'd700, -32'd3746},
{-32'd1966, -32'd12438, 32'd7231, 32'd2569},
{-32'd6440, -32'd9260, 32'd7675, -32'd424},
{32'd8551, 32'd1194, -32'd2227, 32'd320},
{32'd7522, 32'd4273, -32'd4136, -32'd2240},
{-32'd2478, -32'd15529, 32'd2060, 32'd11321},
{32'd3965, -32'd5781, -32'd9173, -32'd1665},
{-32'd6307, 32'd17277, 32'd4184, -32'd800},
{32'd6622, -32'd8554, 32'd6397, 32'd7430},
{-32'd10591, -32'd9737, 32'd25, -32'd2729},
{-32'd5816, 32'd3050, -32'd3727, -32'd1016},
{32'd13184, 32'd8157, -32'd1417, -32'd1862},
{32'd18366, -32'd9596, 32'd1733, -32'd93},
{-32'd4142, -32'd697, -32'd6703, 32'd65},
{-32'd9304, -32'd10593, -32'd11134, -32'd1387},
{-32'd9920, 32'd6549, -32'd1056, 32'd931},
{32'd5073, -32'd2941, -32'd7059, 32'd1176},
{32'd5112, -32'd11836, 32'd2225, 32'd2396},
{32'd12612, -32'd3929, -32'd9301, -32'd2107},
{32'd14701, -32'd114, 32'd8624, -32'd6367},
{32'd19927, -32'd4043, 32'd1285, -32'd415},
{-32'd223, -32'd2732, -32'd1566, -32'd3396},
{32'd12200, 32'd4727, 32'd7328, -32'd1031},
{-32'd23740, -32'd4329, -32'd8461, 32'd6537},
{-32'd16955, -32'd1244, -32'd1186, -32'd3569},
{-32'd15502, 32'd3175, 32'd1670, 32'd7586},
{32'd7411, 32'd9601, -32'd3542, -32'd9807},
{32'd8273, 32'd107, 32'd419, 32'd1304},
{-32'd4122, 32'd216, 32'd3126, 32'd4805},
{32'd11070, 32'd6684, 32'd3830, 32'd3550},
{32'd3246, 32'd1496, 32'd8809, -32'd5342},
{32'd8163, -32'd8188, -32'd14929, -32'd3978},
{-32'd5929, -32'd2185, -32'd591, -32'd775},
{-32'd2686, 32'd255, 32'd4423, 32'd2240},
{32'd6782, 32'd246, 32'd2827, 32'd5555},
{32'd1723, -32'd6786, 32'd3827, 32'd3310},
{32'd645, -32'd9696, -32'd2907, -32'd5476},
{-32'd7542, -32'd3175, 32'd1092, 32'd1022},
{32'd8191, -32'd1476, -32'd6922, -32'd7775},
{-32'd8636, -32'd332, -32'd2363, 32'd8325},
{32'd3969, 32'd7919, -32'd2719, -32'd9852},
{-32'd3008, -32'd7632, -32'd4584, -32'd4781},
{32'd4289, -32'd1054, -32'd1079, 32'd1553},
{32'd5749, -32'd6470, -32'd2951, -32'd346},
{32'd2544, -32'd2827, -32'd942, -32'd4007},
{32'd11569, -32'd5265, -32'd13640, 32'd3269},
{32'd2402, 32'd101, 32'd2595, 32'd9583},
{32'd1714, 32'd2004, -32'd1114, 32'd87},
{-32'd4351, 32'd6860, 32'd3713, -32'd5600},
{32'd9229, 32'd4312, -32'd4889, 32'd345},
{32'd9198, -32'd5670, -32'd6930, 32'd618},
{-32'd7675, -32'd4733, -32'd4891, -32'd5451},
{-32'd18935, 32'd6044, 32'd4008, -32'd1462},
{32'd7732, -32'd13568, 32'd11282, 32'd4968},
{-32'd12990, 32'd2490, 32'd7392, -32'd1035},
{-32'd10920, 32'd1332, -32'd841, 32'd2928},
{32'd10498, -32'd4256, -32'd482, 32'd404},
{-32'd1693, -32'd1578, 32'd3901, -32'd1308},
{32'd333, 32'd17833, -32'd8534, -32'd4978},
{32'd7795, -32'd8477, 32'd7135, -32'd6775},
{32'd16940, -32'd1875, 32'd7429, 32'd367},
{-32'd1666, -32'd1571, -32'd270, -32'd5333},
{-32'd7892, -32'd14294, -32'd2075, 32'd1983},
{32'd2265, 32'd8391, -32'd11858, -32'd8352},
{-32'd2233, -32'd3318, 32'd5249, 32'd1260},
{-32'd13122, 32'd1907, -32'd2052, 32'd1806},
{32'd115, -32'd541, -32'd6243, 32'd28},
{-32'd16307, -32'd11831, 32'd3486, 32'd339},
{32'd1127, 32'd9908, 32'd4206, 32'd6763},
{-32'd18938, -32'd6758, -32'd6308, -32'd4959},
{32'd15432, 32'd9782, 32'd7656, 32'd1804},
{-32'd1702, -32'd11845, -32'd3656, 32'd2568},
{32'd6925, -32'd785, 32'd14020, -32'd1335},
{32'd490, 32'd13018, -32'd2894, 32'd81},
{32'd9849, 32'd5053, -32'd2630, -32'd3253},
{-32'd3048, -32'd3726, -32'd7748, 32'd3414},
{32'd10211, -32'd1250, -32'd1025, 32'd1992},
{32'd5062, -32'd6903, -32'd2875, -32'd219},
{-32'd2830, 32'd2165, -32'd4235, -32'd547},
{-32'd6226, 32'd918, -32'd5679, 32'd5112},
{-32'd6063, 32'd4299, 32'd1556, 32'd1115},
{32'd7178, 32'd7570, 32'd7220, 32'd11108},
{-32'd5083, 32'd1806, -32'd5694, -32'd1555},
{-32'd2875, -32'd4738, 32'd3645, -32'd3940},
{32'd2466, -32'd15911, 32'd3064, 32'd138},
{32'd6301, 32'd6994, 32'd1846, 32'd2052},
{32'd8845, 32'd7992, 32'd833, 32'd5601},
{-32'd3623, -32'd121, -32'd3910, 32'd3101},
{32'd230, -32'd3541, -32'd540, -32'd5844},
{32'd7128, -32'd13600, -32'd7599, -32'd2244},
{32'd9184, -32'd170, -32'd3278, 32'd3136},
{-32'd2026, 32'd4636, -32'd5293, 32'd3173},
{32'd4423, -32'd7123, 32'd6769, 32'd7337},
{32'd159, -32'd7718, 32'd4262, 32'd3667},
{32'd1724, -32'd7156, 32'd10076, 32'd1969},
{32'd6762, 32'd5055, -32'd845, -32'd2138},
{-32'd5455, -32'd545, 32'd1799, -32'd312},
{-32'd8644, -32'd10007, -32'd5460, -32'd1863},
{-32'd6792, 32'd9693, 32'd481, -32'd8435},
{-32'd421, -32'd2786, 32'd3594, 32'd226},
{32'd12122, 32'd10943, -32'd8750, -32'd6991},
{32'd7598, 32'd10321, -32'd2771, -32'd1552},
{-32'd10427, 32'd3467, -32'd2514, -32'd3181},
{32'd5962, -32'd2527, -32'd1479, 32'd8559},
{32'd1565, -32'd1738, -32'd4714, 32'd2765},
{32'd8077, 32'd4507, 32'd596, -32'd3967},
{32'd12502, -32'd4595, -32'd597, -32'd1207},
{-32'd12906, -32'd2861, 32'd5807, 32'd429},
{32'd1438, -32'd4175, 32'd750, 32'd10882},
{-32'd9309, 32'd2637, -32'd1416, -32'd7085},
{32'd1497, -32'd3900, -32'd4302, -32'd1754},
{32'd5410, -32'd1128, 32'd2310, -32'd445},
{-32'd2493, 32'd2535, -32'd1774, 32'd3286},
{32'd8548, -32'd6070, -32'd1155, -32'd2029},
{-32'd8262, 32'd3496, -32'd2470, 32'd5841},
{-32'd5060, -32'd11199, 32'd6526, 32'd5946},
{-32'd7787, -32'd3508, -32'd2859, -32'd5641},
{-32'd662, 32'd821, 32'd4443, 32'd2603},
{32'd17596, 32'd4397, -32'd5011, -32'd5259},
{-32'd1246, 32'd7547, 32'd9691, -32'd3795},
{-32'd187, -32'd4062, 32'd6627, 32'd6305},
{-32'd3438, 32'd9262, 32'd3918, -32'd2308},
{32'd6547, -32'd3326, 32'd2691, -32'd2511},
{-32'd5133, 32'd1062, 32'd3112, 32'd65},
{32'd1017, -32'd3402, -32'd6695, -32'd2360},
{-32'd9117, -32'd1312, -32'd1444, 32'd1144},
{32'd7313, 32'd1549, -32'd8767, -32'd7065},
{32'd10539, -32'd18131, -32'd1930, 32'd8606},
{32'd3812, 32'd4548, -32'd4805, -32'd1420},
{-32'd13415, -32'd4629, 32'd800, -32'd6250},
{-32'd2721, 32'd8379, 32'd1617, 32'd1349},
{-32'd3211, 32'd13364, 32'd6132, 32'd3308},
{-32'd8969, 32'd5298, -32'd1711, 32'd2683},
{-32'd2603, -32'd1367, -32'd7516, 32'd4544},
{32'd82, 32'd8718, -32'd2747, -32'd105},
{32'd1118, -32'd216, -32'd4739, -32'd11332},
{32'd19307, 32'd771, -32'd5885, -32'd863},
{32'd9649, 32'd9756, -32'd7586, 32'd1375},
{32'd3611, -32'd577, 32'd321, -32'd3719},
{-32'd8697, -32'd14468, 32'd1564, -32'd5999},
{32'd709, -32'd4002, -32'd5309, 32'd3489},
{32'd1390, 32'd11373, -32'd969, -32'd1997},
{-32'd1706, -32'd1333, 32'd6967, -32'd1609},
{-32'd5082, -32'd718, 32'd1973, -32'd6000},
{-32'd6823, 32'd2768, -32'd2585, -32'd432},
{-32'd683, -32'd11205, 32'd455, 32'd1709},
{-32'd9977, -32'd5772, 32'd9600, -32'd2709},
{32'd11230, 32'd1628, 32'd1178, -32'd636},
{32'd10698, -32'd5924, -32'd12101, -32'd944},
{-32'd8788, 32'd7100, -32'd3355, 32'd1581},
{-32'd5215, -32'd14394, 32'd2799, -32'd1907},
{32'd4293, -32'd5055, -32'd7975, -32'd5700},
{-32'd10957, -32'd1945, 32'd6430, 32'd3449},
{32'd8914, 32'd2517, 32'd11379, 32'd9551},
{32'd5304, 32'd111, 32'd3170, 32'd4789},
{-32'd14549, 32'd1881, -32'd5151, 32'd638},
{-32'd5604, -32'd3291, -32'd3752, 32'd11707},
{-32'd13688, -32'd3740, -32'd2968, 32'd5136},
{-32'd12867, -32'd746, 32'd1582, 32'd1667},
{-32'd6934, -32'd13743, 32'd3309, -32'd3150},
{-32'd701, 32'd9461, 32'd122, 32'd2126},
{32'd7917, 32'd9728, 32'd1649, 32'd5977},
{-32'd12703, -32'd6333, 32'd4701, -32'd525},
{-32'd7323, -32'd6826, -32'd256, -32'd369},
{32'd3433, -32'd294, -32'd3857, 32'd1555},
{32'd3891, 32'd1735, -32'd24, 32'd1443},
{32'd23647, -32'd5214, 32'd13972, 32'd7015},
{32'd4595, -32'd2565, -32'd4600, -32'd5172},
{-32'd21, -32'd13160, -32'd1947, 32'd7359},
{-32'd16123, -32'd1217, 32'd2420, 32'd8171},
{-32'd1605, 32'd8824, 32'd4902, 32'd5976},
{-32'd8171, 32'd2977, 32'd4855, 32'd2061},
{32'd4561, -32'd5211, 32'd3295, 32'd7266},
{-32'd689, -32'd288, -32'd148, -32'd1753},
{-32'd4116, 32'd2264, 32'd7774, 32'd5306},
{32'd859, 32'd7225, -32'd2404, -32'd3195},
{32'd572, -32'd5355, 32'd1722, -32'd9197},
{32'd3432, 32'd7478, 32'd4185, -32'd6145},
{-32'd11586, -32'd4660, -32'd1593, -32'd4426},
{-32'd8305, 32'd1020, 32'd3078, -32'd2890},
{-32'd2344, -32'd2296, -32'd4360, 32'd1080},
{32'd1931, 32'd4899, -32'd1648, -32'd1188},
{-32'd1819, -32'd12055, -32'd6458, 32'd5111},
{-32'd6463, -32'd10889, 32'd6506, -32'd206},
{32'd7663, 32'd27452, -32'd2035, -32'd3829},
{32'd6743, 32'd2260, 32'd5255, 32'd10004},
{-32'd3914, -32'd2727, -32'd998, 32'd3636},
{32'd526, -32'd144, -32'd4536, -32'd8330},
{32'd2088, 32'd975, -32'd12809, -32'd2008},
{32'd15274, 32'd3237, -32'd1689, 32'd5846},
{-32'd7867, 32'd4720, -32'd7657, 32'd3745},
{-32'd33, 32'd3440, 32'd6115, 32'd1287},
{-32'd10152, -32'd336, -32'd3720, 32'd1504},
{32'd12369, -32'd4571, 32'd5307, 32'd3361},
{-32'd4903, 32'd9411, 32'd2400, -32'd10779},
{32'd2025, -32'd13364, 32'd243, 32'd961},
{-32'd8688, 32'd505, 32'd2715, 32'd245},
{-32'd8407, -32'd3815, -32'd5627, 32'd5941},
{32'd7918, -32'd4254, -32'd60, -32'd4360},
{-32'd8301, 32'd6759, 32'd8886, 32'd62},
{-32'd1485, 32'd3433, 32'd3686, 32'd7550},
{32'd3261, 32'd3898, -32'd3273, 32'd5513},
{32'd4061, 32'd3241, -32'd689, 32'd5010},
{-32'd12465, 32'd6530, 32'd957, -32'd1317},
{-32'd2051, -32'd4181, 32'd2372, -32'd3083},
{-32'd9382, -32'd1916, 32'd7068, -32'd8569},
{32'd2096, -32'd4086, 32'd5848, 32'd2614},
{32'd10845, 32'd9367, -32'd2856, 32'd1664},
{-32'd10610, 32'd1291, 32'd4689, -32'd2791}
},
{{-32'd3290, 32'd4805, 32'd877, -32'd11126},
{-32'd1437, -32'd13496, -32'd17181, 32'd1679},
{32'd2171, -32'd187, 32'd5308, -32'd4119},
{-32'd3213, 32'd1313, -32'd1242, 32'd1418},
{32'd12008, 32'd1828, 32'd8541, 32'd8200},
{-32'd5590, -32'd12175, -32'd2544, 32'd4764},
{32'd10740, 32'd9266, 32'd6635, -32'd5182},
{-32'd21519, 32'd8932, 32'd1760, -32'd8887},
{32'd3631, 32'd2084, 32'd8491, -32'd1107},
{32'd15208, 32'd5446, 32'd4822, 32'd8405},
{-32'd2366, -32'd464, -32'd2448, 32'd3857},
{32'd904, -32'd7445, -32'd12324, 32'd590},
{-32'd6094, -32'd7032, 32'd19483, 32'd10048},
{32'd8830, -32'd3177, 32'd6185, 32'd5902},
{32'd3282, 32'd438, 32'd6793, 32'd4998},
{-32'd3930, 32'd1688, 32'd562, 32'd8917},
{32'd13677, -32'd8534, 32'd13082, -32'd2517},
{-32'd9790, 32'd10824, 32'd7372, 32'd459},
{32'd972, -32'd8018, 32'd11030, -32'd1179},
{32'd1009, -32'd3733, 32'd5940, -32'd5434},
{-32'd8243, -32'd514, -32'd17053, 32'd3578},
{-32'd10160, -32'd10070, -32'd9381, -32'd9086},
{-32'd19187, -32'd4831, -32'd4243, 32'd792},
{-32'd12329, 32'd4596, 32'd3263, -32'd6092},
{32'd5200, -32'd686, -32'd1531, 32'd11676},
{-32'd3363, -32'd6449, -32'd338, -32'd10200},
{-32'd15946, -32'd2213, -32'd8002, -32'd8543},
{-32'd75, 32'd11191, -32'd2208, 32'd1913},
{32'd5211, -32'd13933, 32'd4365, -32'd3748},
{-32'd8391, -32'd11489, -32'd5268, -32'd4846},
{32'd8709, -32'd7278, 32'd5418, 32'd2342},
{-32'd7360, 32'd6972, -32'd14312, -32'd7858},
{32'd12019, -32'd1323, -32'd734, -32'd8122},
{-32'd6848, -32'd1049, 32'd7493, 32'd4757},
{32'd2794, 32'd4188, 32'd5123, 32'd8497},
{32'd2168, -32'd4329, 32'd526, 32'd31},
{32'd9436, 32'd5300, 32'd10270, -32'd2696},
{32'd16931, 32'd5081, -32'd1776, -32'd745},
{32'd8450, 32'd2259, 32'd8114, -32'd2190},
{-32'd3471, 32'd6782, 32'd2597, -32'd3985},
{-32'd3860, -32'd5809, 32'd2501, 32'd2471},
{-32'd11406, 32'd7559, 32'd8275, 32'd8449},
{32'd11472, -32'd9105, -32'd2637, 32'd2546},
{-32'd11735, -32'd1973, -32'd163, 32'd9354},
{-32'd8732, -32'd9769, -32'd700, -32'd6875},
{32'd2737, -32'd2395, -32'd1858, 32'd12110},
{-32'd16407, -32'd2195, 32'd7340, -32'd6504},
{-32'd15162, 32'd1897, 32'd1893, -32'd1552},
{32'd22097, -32'd98, 32'd11630, 32'd1155},
{-32'd1563, -32'd800, -32'd6753, 32'd2205},
{-32'd1233, -32'd98, 32'd10635, -32'd190},
{32'd7028, -32'd5528, -32'd12549, -32'd2686},
{-32'd7651, -32'd893, -32'd6226, 32'd3707},
{32'd1178, 32'd2952, -32'd1384, -32'd4187},
{-32'd15409, -32'd8210, 32'd4633, 32'd13168},
{32'd2837, -32'd7539, -32'd3371, -32'd6635},
{32'd13879, 32'd3092, 32'd19643, 32'd3479},
{-32'd2491, -32'd4224, 32'd725, -32'd16153},
{-32'd7692, 32'd154, -32'd13512, 32'd747},
{32'd4571, -32'd930, -32'd6700, 32'd6563},
{-32'd12556, -32'd2416, -32'd7859, -32'd2397},
{-32'd6727, 32'd5959, 32'd5363, 32'd11601},
{32'd2618, -32'd6389, 32'd3785, -32'd3624},
{32'd3237, 32'd4938, 32'd5472, 32'd2109},
{32'd1160, 32'd1127, 32'd3536, 32'd10478},
{32'd4618, 32'd2149, 32'd7126, 32'd2865},
{-32'd6873, -32'd10109, 32'd857, -32'd227},
{-32'd3116, -32'd3350, -32'd7755, 32'd2573},
{-32'd6184, 32'd3820, -32'd6263, -32'd13037},
{-32'd4934, -32'd8505, 32'd7561, -32'd2527},
{-32'd16634, -32'd431, -32'd5477, -32'd1443},
{-32'd4990, -32'd4739, -32'd12760, 32'd1206},
{-32'd12809, 32'd6170, -32'd8183, 32'd6292},
{32'd2805, 32'd2228, 32'd131, 32'd7091},
{32'd8009, -32'd3709, -32'd8200, -32'd10515},
{-32'd7867, -32'd7569, -32'd1554, -32'd7312},
{-32'd14457, -32'd7248, 32'd1075, 32'd3322},
{-32'd3625, -32'd6947, 32'd8835, -32'd6537},
{32'd10304, 32'd4840, 32'd12951, 32'd6021},
{32'd7122, 32'd9272, -32'd6579, 32'd1031},
{32'd5951, 32'd16055, 32'd13185, -32'd2053},
{-32'd1082, 32'd7991, 32'd6635, 32'd4665},
{32'd8115, -32'd10291, -32'd13355, -32'd2884},
{32'd3932, 32'd1103, -32'd1334, 32'd11412},
{-32'd5763, -32'd4255, -32'd23399, 32'd897},
{32'd2260, 32'd2331, -32'd2493, 32'd10076},
{32'd13047, -32'd9195, 32'd22523, -32'd2932},
{-32'd3269, -32'd7402, 32'd5747, -32'd11012},
{-32'd5707, -32'd3305, 32'd10350, -32'd5896},
{-32'd10321, -32'd8110, -32'd3580, -32'd12532},
{32'd12834, -32'd13471, 32'd9718, 32'd5803},
{32'd920, 32'd1567, 32'd6027, 32'd10937},
{32'd4448, 32'd2130, 32'd3154, 32'd7367},
{32'd6174, -32'd5360, 32'd2750, 32'd16309},
{-32'd9208, 32'd3796, 32'd327, 32'd3022},
{-32'd5990, -32'd7040, -32'd682, -32'd2949},
{32'd11239, 32'd1414, 32'd8928, -32'd3187},
{-32'd14860, -32'd15914, -32'd4054, -32'd8819},
{32'd5678, 32'd7959, -32'd2379, -32'd2878},
{32'd7818, 32'd1670, 32'd7199, -32'd3466},
{-32'd6182, -32'd5213, -32'd9610, -32'd1879},
{-32'd10189, -32'd9656, -32'd3762, 32'd15432},
{-32'd5645, -32'd3941, 32'd10058, 32'd108},
{32'd10494, 32'd8646, 32'd1877, 32'd13315},
{32'd9040, -32'd4337, -32'd4705, 32'd6005},
{-32'd8376, -32'd12233, -32'd7054, 32'd8564},
{-32'd14286, -32'd12089, 32'd10352, 32'd9245},
{-32'd15597, 32'd13851, 32'd7879, 32'd5878},
{-32'd8871, 32'd1786, 32'd5352, 32'd13267},
{-32'd10374, -32'd6142, -32'd516, -32'd354},
{-32'd6071, -32'd7075, -32'd3857, -32'd455},
{-32'd100, 32'd15, -32'd7661, -32'd1973},
{32'd9565, -32'd952, 32'd6133, 32'd3266},
{32'd6563, 32'd9662, 32'd831, -32'd4410},
{-32'd9991, -32'd7014, 32'd6047, 32'd7320},
{-32'd4324, -32'd233, 32'd965, -32'd966},
{-32'd8071, -32'd9854, -32'd15162, 32'd665},
{32'd13064, -32'd6797, -32'd2474, -32'd3841},
{-32'd8922, 32'd205, 32'd4906, 32'd7327},
{32'd7220, 32'd14996, 32'd1250, 32'd6094},
{-32'd2317, 32'd10256, -32'd2565, -32'd762},
{32'd11356, 32'd4787, 32'd13358, -32'd7214},
{32'd7095, -32'd4813, -32'd18492, -32'd567},
{-32'd3185, -32'd5460, 32'd1279, -32'd10823},
{-32'd12279, -32'd2587, -32'd5011, -32'd4595},
{-32'd2715, 32'd2421, 32'd11185, 32'd2877},
{-32'd5496, -32'd8157, 32'd834, 32'd5249},
{-32'd2608, -32'd3438, -32'd5566, -32'd9184},
{-32'd3964, 32'd2693, 32'd10927, 32'd745},
{-32'd4203, -32'd2171, -32'd5370, 32'd163},
{-32'd7972, 32'd1534, -32'd5977, -32'd2743},
{-32'd13611, -32'd1997, -32'd6726, -32'd3031},
{32'd106, 32'd5296, 32'd762, 32'd9309},
{32'd9433, 32'd11061, -32'd4848, 32'd87},
{32'd4297, -32'd223, -32'd3781, -32'd3385},
{32'd3177, 32'd4519, -32'd7666, -32'd9268},
{-32'd852, -32'd164, 32'd3163, -32'd303},
{32'd4445, -32'd14086, 32'd12593, 32'd181},
{-32'd6376, 32'd941, 32'd5658, -32'd5106},
{-32'd13154, -32'd8672, 32'd1649, 32'd6543},
{32'd10357, 32'd8881, 32'd316, -32'd3962},
{-32'd19641, -32'd15975, 32'd6855, -32'd20708},
{32'd6959, 32'd2790, -32'd8007, 32'd7212},
{-32'd3803, -32'd5628, -32'd8075, 32'd9960},
{32'd77, 32'd7661, 32'd8694, 32'd13542},
{32'd8721, 32'd1106, 32'd5367, 32'd2805},
{-32'd6528, -32'd8307, 32'd2843, 32'd6488},
{32'd2036, 32'd8718, -32'd2781, -32'd6522},
{32'd8953, 32'd3939, 32'd4081, -32'd2259},
{32'd4152, -32'd14595, -32'd8423, -32'd6699},
{-32'd6495, -32'd292, 32'd19326, -32'd2271},
{32'd12136, -32'd3298, 32'd4115, -32'd6387},
{32'd15270, 32'd6373, 32'd7856, 32'd3266},
{32'd6105, -32'd2769, 32'd4290, 32'd4687},
{-32'd5472, -32'd7995, -32'd6357, -32'd7168},
{-32'd4847, -32'd119, 32'd8960, -32'd481},
{32'd6399, 32'd14949, -32'd6741, 32'd3187},
{-32'd3695, 32'd4634, -32'd22812, 32'd6525},
{32'd1673, 32'd6797, 32'd2310, -32'd3489},
{32'd10343, -32'd5753, 32'd1379, -32'd7008},
{-32'd337, 32'd11184, -32'd4682, -32'd6394},
{-32'd623, -32'd13297, 32'd6999, -32'd7397},
{-32'd3968, -32'd8077, 32'd8908, -32'd1206},
{32'd6139, -32'd5231, -32'd9021, -32'd6498},
{-32'd2998, 32'd11024, -32'd8627, 32'd22317},
{32'd5965, 32'd398, -32'd8297, -32'd718},
{-32'd2762, -32'd6900, -32'd5313, 32'd15461},
{-32'd5296, -32'd9690, -32'd8027, -32'd5794},
{-32'd13644, -32'd7669, 32'd4767, 32'd6165},
{-32'd4912, -32'd21, -32'd932, 32'd4568},
{-32'd2503, 32'd4190, -32'd460, 32'd1974},
{32'd1045, 32'd7923, 32'd3115, 32'd1536},
{32'd5096, 32'd11161, 32'd2312, 32'd4786},
{-32'd795, 32'd7248, 32'd5656, -32'd2107},
{32'd7980, 32'd5158, 32'd1529, -32'd11981},
{32'd3028, -32'd8675, 32'd3227, 32'd14964},
{32'd15089, 32'd9529, 32'd6747, 32'd1986},
{-32'd1984, -32'd2922, 32'd570, -32'd18525},
{32'd6580, 32'd4994, -32'd2239, -32'd5157},
{-32'd3725, -32'd14835, 32'd1511, -32'd3873},
{-32'd22488, -32'd7832, -32'd7827, -32'd5184},
{32'd4970, -32'd371, -32'd8520, -32'd483},
{-32'd495, -32'd17789, -32'd19657, -32'd3743},
{32'd4316, -32'd2062, 32'd24142, -32'd3886},
{-32'd12631, -32'd2487, 32'd1084, 32'd12386},
{32'd10544, 32'd2429, 32'd2272, 32'd2444},
{-32'd3498, 32'd5432, -32'd13027, -32'd988},
{32'd2033, -32'd9277, -32'd3473, 32'd11427},
{32'd2545, 32'd3243, 32'd314, -32'd7169},
{-32'd17449, -32'd12981, 32'd1044, -32'd11090},
{-32'd9244, -32'd4277, -32'd472, -32'd768},
{-32'd9919, -32'd6797, 32'd35, -32'd1414},
{-32'd14972, 32'd2777, -32'd10092, 32'd14100},
{32'd20850, 32'd2676, 32'd2508, 32'd7006},
{-32'd3029, -32'd6035, -32'd8533, -32'd6734},
{32'd3850, 32'd1746, -32'd3707, -32'd1539},
{32'd1917, 32'd6374, -32'd4979, 32'd8087},
{32'd4251, -32'd1620, 32'd1151, 32'd8574},
{-32'd17874, 32'd10483, 32'd6737, -32'd7814},
{-32'd7357, -32'd3621, 32'd9887, -32'd1646},
{-32'd2973, -32'd14619, -32'd5182, -32'd6783},
{32'd4235, -32'd1928, -32'd7539, -32'd3978},
{32'd15831, -32'd1986, 32'd5042, -32'd10425},
{32'd6695, 32'd8905, 32'd1650, -32'd2869},
{-32'd15509, -32'd16480, -32'd5950, -32'd8929},
{32'd8212, -32'd7452, -32'd8590, -32'd5462},
{32'd9177, -32'd14865, -32'd11667, 32'd7663},
{-32'd3857, 32'd2034, 32'd5773, -32'd2110},
{-32'd8915, -32'd6208, 32'd11311, -32'd5890},
{32'd11166, -32'd12528, -32'd2980, 32'd4849},
{32'd1262, -32'd1566, 32'd9354, 32'd11704},
{-32'd12068, -32'd1634, 32'd12014, 32'd13504},
{32'd9892, -32'd3132, -32'd5915, -32'd7586},
{-32'd8077, 32'd4826, -32'd7759, -32'd16189},
{-32'd962, -32'd320, 32'd8577, -32'd1185},
{32'd1160, -32'd10693, -32'd2237, 32'd7190},
{32'd7819, 32'd8581, -32'd4300, -32'd12399},
{-32'd12045, 32'd3346, -32'd12978, 32'd3523},
{32'd11800, 32'd1000, 32'd11605, -32'd2551},
{-32'd16482, -32'd4959, -32'd7198, -32'd13421},
{32'd1834, -32'd13947, 32'd5853, -32'd11583},
{32'd1275, 32'd5121, 32'd1169, -32'd11497},
{32'd19, 32'd5560, 32'd13428, -32'd11147},
{32'd1856, 32'd3731, 32'd2524, -32'd4371},
{-32'd4978, -32'd12072, -32'd4270, 32'd14666},
{32'd8642, -32'd7638, 32'd7471, 32'd1323},
{32'd731, -32'd13544, 32'd3163, -32'd12673},
{-32'd4153, 32'd11535, -32'd5663, 32'd10257},
{-32'd13463, -32'd4806, 32'd7768, 32'd3144},
{32'd9262, 32'd2040, -32'd646, 32'd1324},
{-32'd10458, 32'd3503, -32'd5159, -32'd3486},
{32'd15356, 32'd14089, 32'd4202, 32'd11610},
{-32'd843, 32'd3348, 32'd4317, -32'd6556},
{32'd1791, -32'd918, -32'd14120, 32'd1502},
{-32'd2093, -32'd7592, -32'd780, -32'd5797},
{32'd1900, -32'd8066, -32'd3464, -32'd8013},
{-32'd8817, 32'd587, -32'd2517, 32'd7339},
{32'd8375, 32'd2549, 32'd5435, 32'd8569},
{32'd244, -32'd4083, -32'd10406, -32'd5074},
{32'd1175, -32'd8129, -32'd40, 32'd516},
{-32'd2454, -32'd1610, 32'd1459, 32'd2878},
{32'd5482, -32'd6093, 32'd10603, -32'd11090},
{-32'd5150, -32'd11444, -32'd2650, 32'd3327},
{32'd9583, -32'd13414, 32'd15989, 32'd15331},
{32'd9158, 32'd6574, 32'd8565, 32'd6304},
{32'd316, 32'd8660, -32'd677, -32'd13440},
{-32'd5543, -32'd1322, -32'd1937, -32'd3364},
{-32'd6069, -32'd13466, -32'd12553, -32'd4731},
{-32'd11389, -32'd8829, -32'd4844, 32'd54},
{32'd846, 32'd3581, 32'd13887, 32'd4277},
{-32'd10327, 32'd3369, 32'd1654, 32'd7105},
{-32'd1787, 32'd3519, -32'd3338, 32'd0},
{-32'd80, 32'd3226, -32'd4903, -32'd6901},
{-32'd3999, 32'd6331, 32'd13399, -32'd629},
{-32'd837, -32'd3656, 32'd3503, 32'd1665},
{32'd2984, 32'd1703, 32'd5028, -32'd1305},
{32'd6751, 32'd4552, 32'd3810, 32'd15902},
{32'd3951, -32'd3319, 32'd2367, 32'd2352},
{-32'd9309, -32'd9697, -32'd10, 32'd535},
{32'd6695, 32'd6784, -32'd3271, -32'd6221},
{32'd1605, 32'd8341, -32'd1400, 32'd8471},
{-32'd20473, 32'd442, 32'd1704, 32'd4132},
{32'd11602, 32'd3359, 32'd10247, -32'd4437},
{-32'd14879, 32'd734, 32'd9791, -32'd5752},
{32'd1271, 32'd2174, 32'd839, 32'd2742},
{-32'd688, -32'd4137, -32'd347, -32'd3376},
{-32'd1008, 32'd8769, 32'd2024, -32'd4372},
{32'd6360, 32'd4160, 32'd449, -32'd1033},
{-32'd4362, -32'd5939, -32'd4490, 32'd12694},
{32'd1613, 32'd11897, 32'd4098, -32'd15360},
{-32'd5763, -32'd2002, -32'd7509, -32'd4216},
{32'd2688, 32'd10324, -32'd4496, -32'd5784},
{32'd5496, -32'd19934, 32'd9838, -32'd9544},
{32'd3436, -32'd11612, -32'd6440, 32'd2587},
{-32'd8482, -32'd10782, -32'd3927, 32'd4210},
{-32'd8752, -32'd6895, -32'd3276, -32'd16389},
{32'd9057, 32'd9690, 32'd4687, 32'd7078},
{32'd9228, 32'd4015, -32'd4984, 32'd6395},
{32'd2820, -32'd7474, -32'd7197, -32'd4126},
{-32'd3668, -32'd3935, -32'd4073, 32'd8679},
{32'd2048, -32'd3554, -32'd1547, -32'd8316},
{32'd9715, 32'd5633, -32'd3084, 32'd8069},
{-32'd8072, 32'd8368, -32'd1678, -32'd3880},
{32'd2660, 32'd8698, -32'd2559, 32'd9697},
{32'd533, 32'd46, -32'd4304, -32'd776},
{-32'd814, -32'd2296, 32'd6984, -32'd1969},
{-32'd3391, 32'd6598, -32'd5365, -32'd10331},
{-32'd50, 32'd2888, 32'd9904, -32'd3980},
{-32'd5345, 32'd13081, 32'd5844, -32'd8396},
{-32'd2803, 32'd10734, -32'd14138, -32'd7633},
{32'd442, -32'd8495, 32'd13404, 32'd2550},
{32'd7263, 32'd18024, -32'd7407, 32'd3943},
{-32'd691, -32'd14617, 32'd5851, 32'd12985},
{-32'd11130, 32'd3580, -32'd3140, -32'd10938},
{-32'd13618, -32'd1992, 32'd1860, 32'd4035},
{-32'd9888, -32'd5604, 32'd8564, -32'd7284},
{32'd83, -32'd7516, 32'd5022, 32'd10889},
{32'd5361, -32'd3815, -32'd5292, -32'd8173},
{-32'd733, 32'd10515, -32'd1714, 32'd7677},
{-32'd4244, 32'd9189, 32'd6236, -32'd12125}
},
{{32'd9370, 32'd3031, 32'd2261, 32'd2886},
{32'd2679, -32'd1910, 32'd7396, -32'd2463},
{32'd648, -32'd12879, -32'd1637, 32'd5075},
{32'd9477, 32'd2784, -32'd1654, 32'd3577},
{32'd5822, -32'd3955, 32'd495, 32'd3161},
{-32'd1471, -32'd1835, 32'd2759, -32'd4864},
{-32'd6784, -32'd8730, 32'd854, 32'd1316},
{-32'd11622, -32'd5530, 32'd686, -32'd3278},
{32'd2752, -32'd8078, 32'd4104, 32'd2212},
{32'd18186, 32'd3703, 32'd1469, 32'd8766},
{32'd4609, -32'd4548, 32'd6984, -32'd4150},
{-32'd5313, -32'd691, -32'd4519, -32'd4432},
{32'd12670, -32'd8592, -32'd9488, 32'd726},
{-32'd5652, -32'd4499, -32'd4846, 32'd1546},
{-32'd10484, -32'd6678, -32'd6787, -32'd4078},
{32'd694, -32'd3176, -32'd7740, -32'd1288},
{32'd2448, 32'd8329, -32'd369, -32'd1598},
{32'd8566, 32'd3345, -32'd1318, 32'd38},
{32'd6660, -32'd422, -32'd6498, 32'd2558},
{-32'd3695, -32'd86, -32'd7948, 32'd2331},
{32'd3952, -32'd5922, -32'd13610, 32'd4256},
{32'd5742, 32'd239, -32'd12114, -32'd2636},
{-32'd3449, -32'd3260, -32'd8303, -32'd6263},
{32'd4582, 32'd2615, -32'd3185, -32'd6932},
{32'd13602, 32'd1879, -32'd31, 32'd1412},
{-32'd3828, -32'd5578, -32'd1351, -32'd5840},
{-32'd8076, 32'd3952, 32'd6958, -32'd5406},
{32'd11941, 32'd6440, 32'd1476, -32'd5236},
{-32'd4363, 32'd1086, 32'd5107, 32'd1479},
{-32'd12276, -32'd8813, -32'd7540, 32'd5839},
{32'd2101, -32'd5634, -32'd3596, -32'd4796},
{32'd274, -32'd4346, -32'd3283, -32'd5928},
{32'd13186, 32'd1915, 32'd1711, 32'd5907},
{32'd4119, 32'd178, -32'd8468, -32'd3002},
{32'd17530, 32'd4598, 32'd10723, 32'd684},
{-32'd14898, -32'd67, -32'd2196, -32'd2484},
{-32'd16, -32'd1405, -32'd2665, -32'd849},
{32'd7447, -32'd3489, -32'd520, 32'd7028},
{32'd6941, 32'd1062, 32'd193, 32'd510},
{32'd5738, 32'd5260, 32'd2326, -32'd5502},
{32'd1934, 32'd4505, -32'd4908, 32'd2207},
{32'd6442, -32'd6887, 32'd4359, 32'd2702},
{32'd8814, 32'd7347, 32'd2728, 32'd117},
{-32'd4119, -32'd14786, -32'd8979, -32'd1761},
{-32'd16866, -32'd6262, -32'd8145, -32'd982},
{32'd2212, -32'd5542, -32'd5699, 32'd2613},
{32'd11640, 32'd197, -32'd7298, -32'd6118},
{-32'd6463, 32'd6108, 32'd16, -32'd2030},
{-32'd2951, 32'd8751, 32'd3390, 32'd4638},
{-32'd6332, -32'd5668, -32'd3221, 32'd1621},
{-32'd9013, -32'd2717, -32'd3637, -32'd2349},
{32'd3002, -32'd4305, 32'd4057, 32'd1955},
{32'd4522, 32'd4161, -32'd1961, -32'd2919},
{32'd4234, -32'd7961, 32'd306, -32'd729},
{32'd4382, -32'd3032, -32'd1092, -32'd2875},
{-32'd4381, 32'd3965, 32'd6827, -32'd363},
{32'd8842, 32'd2041, 32'd2696, 32'd2130},
{-32'd7253, -32'd4496, -32'd3965, -32'd3581},
{-32'd1935, -32'd4449, -32'd3709, -32'd4995},
{-32'd1215, 32'd7615, 32'd188, -32'd5204},
{-32'd4009, 32'd4962, -32'd98, -32'd4141},
{32'd4015, -32'd827, 32'd6427, -32'd1176},
{-32'd6253, 32'd551, -32'd1614, -32'd8219},
{-32'd2191, -32'd13157, 32'd5966, 32'd767},
{32'd5553, 32'd4933, -32'd6546, 32'd8051},
{32'd2693, -32'd5219, 32'd3684, 32'd3294},
{32'd785, 32'd5279, -32'd2556, -32'd166},
{-32'd8923, -32'd10993, 32'd2948, -32'd2149},
{32'd5016, -32'd6144, -32'd7834, 32'd432},
{-32'd1743, -32'd2190, -32'd1729, -32'd2307},
{32'd5073, -32'd10694, 32'd1375, -32'd2854},
{32'd7798, -32'd8831, 32'd4938, -32'd277},
{-32'd2371, 32'd494, 32'd4779, -32'd2145},
{-32'd4657, 32'd438, 32'd3385, 32'd4988},
{32'd309, -32'd380, 32'd1761, 32'd6551},
{32'd6406, 32'd2919, -32'd9742, 32'd832},
{-32'd668, 32'd1251, -32'd955, -32'd93},
{-32'd6221, 32'd3183, 32'd9517, -32'd6446},
{-32'd390, 32'd258, -32'd4683, 32'd2133},
{32'd63, -32'd650, 32'd2894, -32'd2991},
{32'd1404, -32'd1504, 32'd681, 32'd658},
{-32'd3163, 32'd3775, 32'd769, -32'd1596},
{32'd911, 32'd1808, -32'd611, -32'd4169},
{32'd7859, -32'd7092, 32'd5664, 32'd1214},
{32'd1759, -32'd3359, 32'd1614, -32'd2718},
{-32'd8033, -32'd8162, -32'd1276, -32'd365},
{32'd4182, 32'd2438, 32'd4230, 32'd1979},
{-32'd2399, -32'd10029, 32'd1122, -32'd10550},
{-32'd657, 32'd1805, -32'd3827, -32'd1542},
{-32'd6226, 32'd4808, -32'd4465, 32'd686},
{32'd10896, 32'd819, 32'd6151, 32'd6902},
{32'd289, -32'd1623, -32'd1115, 32'd5725},
{32'd2283, -32'd1141, 32'd164, 32'd8550},
{32'd15068, 32'd11626, 32'd4095, 32'd9834},
{32'd2294, 32'd3875, 32'd2200, -32'd4419},
{32'd6732, 32'd844, -32'd3641, -32'd645},
{32'd5128, 32'd364, 32'd3274, -32'd4486},
{-32'd12068, 32'd2342, -32'd4577, 32'd2413},
{-32'd1485, -32'd4318, 32'd10515, -32'd339},
{32'd7307, -32'd2674, 32'd1014, 32'd4763},
{32'd1873, 32'd19442, -32'd8869, -32'd718},
{32'd4160, -32'd14810, -32'd8071, -32'd6358},
{-32'd2531, 32'd5714, -32'd1154, -32'd2839},
{32'd255, -32'd1772, 32'd11371, 32'd786},
{32'd11453, 32'd7307, 32'd7853, -32'd950},
{32'd3815, -32'd6949, -32'd520, -32'd1689},
{-32'd7776, 32'd3935, 32'd2043, -32'd4832},
{32'd218, -32'd8723, -32'd2078, 32'd3821},
{32'd6810, 32'd9314, 32'd1389, -32'd2062},
{-32'd10407, 32'd4598, -32'd2324, -32'd1705},
{-32'd367, 32'd6272, -32'd3224, -32'd2292},
{32'd7244, 32'd10616, 32'd1111, 32'd1847},
{-32'd885, -32'd3650, 32'd4175, 32'd1538},
{32'd5527, 32'd13656, 32'd4365, 32'd3234},
{32'd2682, -32'd3700, -32'd1721, -32'd7411},
{-32'd3830, 32'd6890, -32'd1928, 32'd3504},
{32'd1993, 32'd2502, 32'd3973, -32'd1545},
{-32'd1055, 32'd5426, 32'd2831, -32'd3689},
{-32'd875, -32'd894, 32'd3783, 32'd1523},
{32'd6555, 32'd7190, 32'd2508, 32'd4683},
{32'd9180, -32'd1420, -32'd876, 32'd702},
{32'd6412, 32'd7875, -32'd7938, -32'd1231},
{32'd4485, -32'd3799, 32'd951, -32'd1619},
{32'd1407, 32'd7287, 32'd1346, -32'd4421},
{32'd5960, 32'd2604, 32'd2790, 32'd1795},
{32'd3152, -32'd2870, -32'd1194, 32'd9877},
{-32'd1466, 32'd987, -32'd9206, -32'd8480},
{-32'd4494, -32'd5542, -32'd2067, -32'd7185},
{32'd9222, 32'd2886, 32'd4061, -32'd4308},
{32'd10192, -32'd11074, 32'd1482, 32'd4120},
{-32'd8964, -32'd2510, 32'd6939, -32'd1678},
{-32'd8308, -32'd13844, 32'd1540, -32'd5422},
{-32'd7363, -32'd6592, 32'd5245, -32'd1770},
{32'd2572, 32'd2672, 32'd366, 32'd1835},
{32'd5885, 32'd1119, -32'd917, -32'd3149},
{32'd2510, 32'd449, -32'd5666, -32'd2728},
{-32'd7021, 32'd6962, -32'd3599, 32'd6830},
{-32'd7195, -32'd12082, 32'd7343, -32'd2749},
{32'd5944, 32'd2817, 32'd3318, 32'd448},
{-32'd4591, 32'd2398, 32'd8815, -32'd765},
{-32'd11129, 32'd353, 32'd3227, -32'd2107},
{-32'd1373, -32'd3337, -32'd2726, -32'd6444},
{32'd7476, -32'd17871, 32'd1831, 32'd4546},
{32'd3755, -32'd4669, 32'd802, 32'd3071},
{32'd15702, 32'd7727, 32'd2900, 32'd2594},
{-32'd1548, 32'd395, 32'd840, 32'd5161},
{-32'd6281, 32'd6993, 32'd4809, -32'd2110},
{32'd6331, -32'd10231, 32'd3868, -32'd503},
{32'd7532, -32'd941, 32'd12158, 32'd5783},
{32'd4147, 32'd879, 32'd5991, -32'd7490},
{-32'd12501, -32'd763, -32'd6845, -32'd2118},
{32'd2458, 32'd1931, -32'd1146, 32'd4978},
{-32'd3305, -32'd275, 32'd5903, 32'd1094},
{32'd4957, -32'd2856, -32'd4205, -32'd577},
{-32'd12257, -32'd8678, -32'd9455, -32'd7428},
{-32'd6046, -32'd11333, 32'd6559, -32'd2766},
{32'd5453, -32'd4335, 32'd5422, -32'd1275},
{-32'd1683, 32'd494, 32'd288, -32'd1502},
{32'd1036, -32'd816, -32'd6558, -32'd2577},
{32'd7314, -32'd1154, 32'd3796, -32'd768},
{-32'd11828, 32'd3791, -32'd1231, -32'd3925},
{32'd1035, 32'd3487, -32'd779, 32'd846},
{-32'd9018, 32'd2726, -32'd1890, -32'd1387},
{-32'd4885, 32'd2339, 32'd4156, -32'd838},
{32'd3642, -32'd9787, 32'd8095, 32'd7950},
{-32'd1873, 32'd1604, -32'd5318, 32'd3726},
{32'd1114, -32'd7375, 32'd13337, 32'd1764},
{-32'd399, -32'd12922, -32'd5485, 32'd2056},
{32'd632, 32'd895, 32'd4993, -32'd856},
{-32'd3534, -32'd4769, 32'd5828, 32'd1721},
{32'd9892, 32'd12930, -32'd3090, -32'd1469},
{-32'd821, 32'd6156, 32'd2415, -32'd1342},
{32'd9914, 32'd1167, 32'd15977, -32'd2234},
{-32'd170, 32'd4025, 32'd4057, -32'd1769},
{32'd5627, -32'd3488, -32'd3238, -32'd2085},
{32'd2644, 32'd993, -32'd3210, 32'd5508},
{-32'd6228, 32'd10887, -32'd1753, 32'd155},
{32'd9978, -32'd9866, -32'd6574, 32'd4004},
{32'd2938, 32'd8232, -32'd1910, -32'd2125},
{-32'd12535, 32'd2501, -32'd7800, -32'd1772},
{-32'd5320, -32'd2573, -32'd4235, -32'd970},
{-32'd1768, -32'd8032, -32'd758, 32'd3740},
{-32'd4446, 32'd1758, -32'd11453, -32'd9817},
{-32'd2107, -32'd1385, -32'd5833, -32'd185},
{32'd3900, -32'd4469, -32'd6502, -32'd3271},
{32'd2140, 32'd314, -32'd522, 32'd2427},
{32'd3802, -32'd4481, -32'd256, 32'd1869},
{-32'd10556, -32'd4964, 32'd2020, -32'd873},
{-32'd2171, 32'd597, 32'd2926, -32'd1681},
{32'd2719, -32'd495, -32'd7641, 32'd4849},
{32'd3316, -32'd718, 32'd1735, -32'd4551},
{-32'd844, -32'd6601, -32'd852, -32'd5326},
{-32'd7156, 32'd3737, 32'd201, -32'd1240},
{32'd3537, -32'd405, 32'd3124, -32'd3298},
{-32'd11349, -32'd10931, 32'd4510, 32'd5304},
{-32'd1465, -32'd4549, -32'd4658, -32'd4667},
{-32'd6210, 32'd5041, 32'd8196, -32'd7528},
{-32'd30, -32'd1267, 32'd817, 32'd8543},
{32'd4481, -32'd7179, -32'd3171, 32'd4012},
{-32'd8573, -32'd6178, -32'd2487, 32'd2534},
{-32'd15708, -32'd324, -32'd7967, -32'd5540},
{32'd7581, 32'd3929, -32'd3342, -32'd800},
{32'd5176, -32'd3641, 32'd4027, -32'd602},
{-32'd4564, 32'd7730, 32'd5991, -32'd3726},
{-32'd4189, 32'd2649, -32'd5197, -32'd4762},
{32'd7157, -32'd1752, 32'd10416, 32'd844},
{32'd1468, 32'd8294, 32'd481, 32'd3773},
{32'd2677, -32'd8829, 32'd1246, -32'd831},
{-32'd2177, 32'd2882, 32'd241, 32'd4379},
{32'd12741, 32'd10556, 32'd9252, -32'd1994},
{32'd869, -32'd1811, -32'd9955, 32'd381},
{-32'd6472, -32'd485, 32'd2199, -32'd362},
{-32'd7030, -32'd8006, -32'd4115, 32'd2993},
{32'd1702, -32'd2022, 32'd8695, 32'd3348},
{-32'd4712, 32'd10124, -32'd4613, -32'd5584},
{32'd4641, -32'd6142, 32'd1027, -32'd3821},
{32'd1473, -32'd1841, 32'd4014, 32'd1891},
{32'd7541, -32'd19646, -32'd1289, -32'd4636},
{-32'd3858, 32'd1634, 32'd11973, 32'd2298},
{-32'd8943, -32'd11014, -32'd14401, -32'd890},
{-32'd8993, 32'd4735, -32'd10871, 32'd362},
{-32'd448, 32'd6256, 32'd13, -32'd952},
{32'd2618, -32'd3888, -32'd3610, 32'd374},
{32'd5045, -32'd5594, -32'd4323, -32'd3690},
{-32'd8592, 32'd1367, -32'd4316, 32'd2645},
{-32'd2026, 32'd171, 32'd5160, 32'd2890},
{-32'd3857, 32'd7988, 32'd4917, 32'd829},
{-32'd15912, -32'd4437, 32'd2361, -32'd5346},
{-32'd3859, 32'd320, -32'd7580, -32'd7655},
{-32'd3597, 32'd124, 32'd3425, 32'd7496},
{32'd5311, -32'd3003, 32'd3679, -32'd6586},
{32'd2375, 32'd5350, 32'd2689, -32'd393},
{32'd6172, -32'd1932, -32'd1356, -32'd1852},
{-32'd11710, 32'd2524, -32'd6744, -32'd5877},
{32'd2981, 32'd535, -32'd7675, -32'd1198},
{32'd290, 32'd6589, -32'd6479, -32'd2604},
{32'd2791, 32'd2390, -32'd1543, -32'd195},
{32'd1882, 32'd6870, -32'd4864, -32'd4940},
{-32'd3591, -32'd6272, 32'd2323, -32'd721},
{-32'd1018, 32'd129, -32'd2046, -32'd3332},
{32'd11919, 32'd465, 32'd4165, -32'd1784},
{-32'd7064, -32'd1153, -32'd3205, -32'd5775},
{-32'd6992, 32'd5784, -32'd9955, -32'd9278},
{32'd2591, 32'd6088, 32'd1144, 32'd7721},
{32'd9971, 32'd7058, 32'd2562, 32'd7350},
{32'd10802, 32'd10358, -32'd50, -32'd3713},
{32'd2506, 32'd4765, 32'd5418, -32'd5394},
{-32'd5723, 32'd8259, 32'd318, 32'd2684},
{32'd2969, 32'd1119, -32'd6305, -32'd3538},
{-32'd3746, -32'd1276, 32'd2203, 32'd3716},
{32'd6522, -32'd3550, 32'd1422, 32'd2641},
{-32'd9629, 32'd7694, -32'd4246, -32'd9872},
{-32'd1475, 32'd9937, -32'd3636, 32'd1587},
{32'd11785, 32'd3222, -32'd7064, 32'd2946},
{-32'd11423, -32'd1152, -32'd4762, 32'd3855},
{32'd3943, 32'd5549, 32'd330, 32'd3021},
{32'd7976, 32'd3167, -32'd4323, 32'd3960},
{-32'd6419, 32'd13252, 32'd3897, 32'd3463},
{32'd3545, 32'd7973, -32'd3308, -32'd6759},
{-32'd3409, 32'd1946, 32'd3036, 32'd4161},
{32'd4221, -32'd3031, 32'd5649, 32'd2310},
{32'd15063, -32'd6893, -32'd7660, -32'd2618},
{-32'd6619, -32'd8870, -32'd2276, 32'd1068},
{-32'd8344, -32'd6051, -32'd4974, -32'd5856},
{-32'd5741, -32'd793, -32'd5724, -32'd1189},
{32'd1309, 32'd1691, -32'd5009, 32'd3790},
{32'd6447, 32'd54, -32'd9612, -32'd3475},
{-32'd249, -32'd7420, -32'd490, -32'd3333},
{32'd698, -32'd10008, -32'd9076, -32'd5703},
{32'd944, 32'd12156, -32'd445, 32'd6332},
{32'd5289, 32'd4367, 32'd6439, -32'd3405},
{-32'd11177, -32'd2056, 32'd13251, 32'd4381},
{-32'd3806, -32'd5364, -32'd5467, 32'd1730},
{-32'd2337, -32'd7722, -32'd4382, -32'd823},
{32'd2790, -32'd7895, -32'd1737, 32'd411},
{-32'd3423, 32'd2853, -32'd10033, 32'd618},
{32'd21461, 32'd4847, 32'd3218, 32'd8988},
{32'd14535, 32'd1739, -32'd537, -32'd427},
{-32'd9625, -32'd1271, -32'd1461, -32'd3260},
{32'd5847, -32'd1004, 32'd5168, -32'd4480},
{32'd8594, 32'd2475, -32'd1810, 32'd923},
{32'd3404, 32'd3357, 32'd6756, 32'd6454},
{32'd9929, -32'd2343, 32'd1782, 32'd8904},
{32'd4914, -32'd4764, 32'd7813, -32'd1215},
{32'd9777, -32'd17880, 32'd4494, 32'd1994},
{-32'd1163, -32'd1915, 32'd3403, -32'd3962},
{32'd10701, 32'd3093, -32'd1571, 32'd714},
{32'd3104, 32'd15487, -32'd5440, -32'd2567},
{32'd2019, 32'd10892, 32'd7782, 32'd295},
{-32'd2478, 32'd8969, -32'd650, -32'd6129},
{32'd2948, -32'd14062, -32'd4922, -32'd2527},
{-32'd8997, 32'd8187, 32'd858, 32'd7718},
{32'd5689, 32'd6109, -32'd2902, -32'd4364},
{32'd6560, -32'd1113, -32'd4723, -32'd1004},
{32'd1060, 32'd2080, 32'd1871, -32'd3765},
{-32'd5093, -32'd5229, 32'd353, -32'd5066},
{32'd4410, -32'd8752, 32'd1264, 32'd37},
{-32'd851, -32'd3278, -32'd3125, 32'd2973},
{32'd3345, -32'd444, 32'd10480, -32'd1968},
{32'd5318, 32'd7134, -32'd7251, -32'd5937}
},
{{-32'd4496, 32'd5105, 32'd618, 32'd4472},
{-32'd9827, -32'd8633, -32'd5870, -32'd5332},
{-32'd1165, -32'd7561, -32'd1050, 32'd323},
{-32'd3406, -32'd4133, 32'd6895, -32'd6952},
{32'd10727, -32'd7543, 32'd4131, 32'd2325},
{-32'd16617, 32'd1444, -32'd8470, -32'd2945},
{32'd9531, -32'd660, 32'd4882, -32'd5116},
{-32'd3107, 32'd5820, -32'd1491, 32'd853},
{32'd9418, 32'd643, 32'd4399, 32'd6418},
{32'd6201, -32'd913, 32'd2974, -32'd1457},
{-32'd6567, 32'd2344, -32'd2145, -32'd3336},
{32'd10002, 32'd2013, -32'd9662, -32'd11549},
{32'd4086, -32'd301, 32'd5219, -32'd7757},
{32'd10129, 32'd10285, -32'd683, 32'd647},
{32'd2803, 32'd5073, -32'd2829, -32'd5180},
{32'd6787, 32'd9786, -32'd5842, 32'd1292},
{-32'd4264, -32'd9416, 32'd5704, -32'd8327},
{-32'd1809, 32'd12474, -32'd6584, 32'd19297},
{32'd12885, 32'd3419, 32'd6479, -32'd11365},
{32'd15219, -32'd11404, -32'd4937, 32'd9795},
{32'd3951, -32'd3779, -32'd6760, -32'd5997},
{-32'd5270, 32'd3554, -32'd912, -32'd948},
{-32'd1797, -32'd7232, 32'd5174, -32'd202},
{-32'd3609, 32'd1685, 32'd8271, 32'd2582},
{32'd5989, 32'd1613, 32'd5327, 32'd620},
{32'd7010, 32'd2636, 32'd10341, -32'd7175},
{-32'd8158, -32'd17538, -32'd5906, 32'd10542},
{-32'd4063, -32'd7402, 32'd65, 32'd3933},
{-32'd2669, -32'd12505, -32'd1055, -32'd7536},
{32'd6335, 32'd3946, 32'd2163, 32'd284},
{32'd9849, 32'd1376, -32'd6540, 32'd8021},
{-32'd874, 32'd1161, 32'd1205, 32'd8113},
{-32'd718, -32'd7695, 32'd1925, -32'd9052},
{32'd2575, -32'd7371, 32'd1119, 32'd3236},
{32'd6457, 32'd3238, 32'd3368, 32'd6694},
{32'd4226, 32'd7124, 32'd6319, 32'd813},
{-32'd6429, -32'd11897, 32'd4309, 32'd7175},
{32'd5309, 32'd2910, 32'd5130, -32'd2160},
{-32'd1407, -32'd9219, -32'd7783, -32'd19563},
{-32'd3078, 32'd9010, -32'd283, 32'd1384},
{-32'd9374, -32'd12983, -32'd5391, 32'd5939},
{32'd6949, 32'd9761, 32'd2169, 32'd6551},
{32'd5621, -32'd1163, -32'd826, -32'd3115},
{32'd11165, 32'd5359, -32'd9451, -32'd5825},
{32'd3164, 32'd8057, 32'd798, -32'd5930},
{32'd9580, -32'd2566, -32'd2906, 32'd597},
{-32'd7050, -32'd1898, 32'd5669, 32'd4717},
{32'd6037, 32'd3832, -32'd4501, 32'd832},
{32'd3061, 32'd6222, -32'd8524, 32'd3878},
{32'd6991, 32'd8274, -32'd4126, 32'd7339},
{32'd4119, -32'd9150, 32'd1018, -32'd1905},
{-32'd538, 32'd623, 32'd642, 32'd13917},
{-32'd4892, -32'd6038, 32'd1556, 32'd1627},
{-32'd4490, -32'd3486, 32'd9926, -32'd5094},
{32'd4535, 32'd10785, -32'd181, 32'd4160},
{-32'd1146, -32'd1698, -32'd6597, -32'd2677},
{-32'd1586, 32'd3029, 32'd5391, -32'd1653},
{-32'd12646, 32'd7026, 32'd1007, -32'd975},
{32'd6903, 32'd5074, -32'd9681, 32'd3555},
{32'd8916, -32'd1288, -32'd817, 32'd7372},
{-32'd4958, 32'd11076, -32'd1074, -32'd881},
{-32'd5541, -32'd3134, -32'd2592, -32'd7773},
{32'd2910, -32'd4030, 32'd3473, -32'd1048},
{32'd13433, -32'd13167, -32'd4272, -32'd6122},
{-32'd11594, -32'd988, -32'd732, 32'd4678},
{32'd5661, 32'd4038, 32'd2573, -32'd3898},
{-32'd800, -32'd12597, -32'd2152, 32'd469},
{-32'd5402, -32'd7724, -32'd935, 32'd12176},
{-32'd13954, -32'd9875, 32'd2281, -32'd1293},
{-32'd3352, -32'd4496, 32'd1009, 32'd10},
{-32'd4748, -32'd8046, -32'd14390, 32'd3989},
{-32'd4077, 32'd2568, 32'd2836, 32'd4521},
{32'd635, -32'd6460, 32'd2742, 32'd11275},
{32'd4208, 32'd1595, 32'd162, -32'd12160},
{-32'd4302, -32'd3133, 32'd9543, -32'd6412},
{-32'd2451, -32'd7876, 32'd2728, -32'd2344},
{-32'd15420, 32'd11805, -32'd2365, 32'd3417},
{32'd4025, 32'd2241, 32'd3562, -32'd10777},
{-32'd1230, 32'd11210, 32'd2734, -32'd8189},
{-32'd1763, 32'd4969, 32'd12836, -32'd1545},
{-32'd7732, -32'd536, -32'd2594, -32'd7185},
{-32'd4326, -32'd6761, 32'd4977, 32'd874},
{32'd4440, -32'd8871, -32'd1139, 32'd1406},
{32'd4460, -32'd3263, -32'd3511, 32'd9372},
{-32'd2697, 32'd9622, 32'd1672, 32'd3207},
{-32'd244, -32'd2347, -32'd1453, -32'd4339},
{32'd14265, -32'd15918, -32'd38, -32'd360},
{-32'd3564, -32'd525, 32'd2284, 32'd2101},
{32'd4941, -32'd7541, -32'd1237, 32'd3047},
{32'd7364, 32'd254, 32'd6646, -32'd9189},
{32'd3660, 32'd7557, -32'd5678, 32'd5140},
{32'd785, 32'd2782, 32'd3342, -32'd7962},
{32'd4902, 32'd8054, 32'd3944, 32'd3072},
{-32'd3366, -32'd950, -32'd12554, 32'd8730},
{-32'd3373, -32'd3020, 32'd4572, 32'd206},
{-32'd1211, -32'd8700, -32'd15703, -32'd4732},
{-32'd3303, -32'd481, 32'd11640, -32'd9036},
{-32'd10485, 32'd8492, -32'd541, 32'd11323},
{-32'd13262, -32'd6215, 32'd1955, 32'd7362},
{32'd4687, 32'd8557, -32'd4872, -32'd10154},
{-32'd9341, 32'd2028, 32'd6949, -32'd2319},
{-32'd3329, 32'd10246, 32'd2530, 32'd10901},
{-32'd5453, -32'd9958, 32'd5110, -32'd304},
{32'd1730, -32'd282, 32'd2634, -32'd12287},
{32'd4083, -32'd511, 32'd9671, 32'd6249},
{32'd7582, 32'd11174, -32'd942, -32'd3752},
{32'd5285, 32'd1624, 32'd5451, 32'd4972},
{32'd877, -32'd10098, -32'd8538, 32'd9282},
{32'd8353, 32'd757, -32'd2693, 32'd4207},
{32'd5499, 32'd869, 32'd5096, -32'd3062},
{-32'd4863, -32'd4452, -32'd5519, 32'd2522},
{-32'd4680, -32'd6081, 32'd6057, -32'd3416},
{32'd10630, -32'd11120, -32'd1408, -32'd5767},
{-32'd4526, -32'd541, 32'd3150, 32'd3296},
{32'd4054, -32'd367, 32'd3996, 32'd2658},
{-32'd9875, -32'd15545, 32'd706, 32'd3756},
{32'd5710, 32'd8840, 32'd10825, 32'd138},
{-32'd2340, 32'd6208, 32'd1001, -32'd139},
{-32'd9939, 32'd7249, -32'd5763, -32'd4110},
{32'd3675, 32'd9447, 32'd2683, 32'd4719},
{32'd6367, -32'd3263, -32'd3510, -32'd4022},
{-32'd2560, 32'd1950, 32'd13055, -32'd7913},
{32'd5898, 32'd1766, 32'd36, 32'd2238},
{32'd112, -32'd12839, 32'd9231, 32'd2105},
{-32'd7925, -32'd5008, -32'd2785, -32'd9534},
{-32'd7478, -32'd8959, -32'd1194, 32'd1025},
{32'd6210, 32'd10476, 32'd5839, 32'd6849},
{32'd1639, -32'd1642, -32'd2992, 32'd2509},
{32'd3711, -32'd11596, -32'd661, -32'd3807},
{-32'd1485, 32'd380, -32'd4149, -32'd1186},
{-32'd3431, 32'd9834, 32'd5432, -32'd4531},
{-32'd9159, 32'd4023, -32'd583, 32'd7182},
{-32'd12300, -32'd3202, -32'd11896, -32'd3967},
{-32'd6033, -32'd15019, -32'd4532, 32'd4260},
{-32'd2743, -32'd9313, 32'd5814, 32'd5976},
{-32'd7974, -32'd1670, 32'd1326, 32'd3342},
{-32'd1626, 32'd11840, 32'd13031, 32'd4736},
{-32'd12202, 32'd1868, 32'd5306, -32'd7538},
{-32'd3173, -32'd4055, -32'd2788, -32'd575},
{-32'd2571, -32'd12286, -32'd7047, 32'd1801},
{32'd7473, -32'd6398, -32'd277, 32'd3928},
{32'd6147, -32'd4607, 32'd191, -32'd3369},
{-32'd2880, 32'd11579, 32'd5295, -32'd6610},
{-32'd3703, 32'd2640, -32'd3329, 32'd4150},
{-32'd3032, 32'd2063, -32'd438, -32'd1812},
{-32'd6622, 32'd3784, -32'd4465, 32'd5629},
{32'd2783, -32'd1509, 32'd2133, 32'd6962},
{32'd8859, -32'd1305, 32'd4181, -32'd4442},
{-32'd4547, -32'd4872, -32'd2653, -32'd1577},
{-32'd11586, 32'd3076, 32'd2196, -32'd4187},
{-32'd5591, -32'd1096, -32'd6508, -32'd651},
{-32'd7193, 32'd2219, 32'd4963, 32'd5769},
{-32'd1917, -32'd925, 32'd3378, -32'd8431},
{32'd354, -32'd7589, -32'd3806, 32'd409},
{-32'd3558, -32'd6410, 32'd1664, -32'd342},
{-32'd3334, -32'd6164, -32'd7426, 32'd1908},
{32'd10373, 32'd11830, 32'd14236, 32'd5260},
{-32'd44, 32'd2736, -32'd3769, 32'd3954},
{-32'd4985, -32'd4306, 32'd4912, -32'd13209},
{32'd6425, 32'd6224, 32'd6294, -32'd3368},
{-32'd5119, 32'd6900, 32'd2945, 32'd4694},
{-32'd5781, -32'd5473, 32'd10551, -32'd5980},
{-32'd4376, -32'd10548, 32'd10486, 32'd17993},
{32'd952, 32'd4643, -32'd18578, -32'd8625},
{32'd7949, 32'd3781, -32'd7497, -32'd3710},
{32'd343, -32'd8320, -32'd4378, -32'd1223},
{32'd9543, 32'd9942, -32'd7808, 32'd3345},
{32'd2844, -32'd970, -32'd10855, -32'd572},
{-32'd3950, -32'd6744, -32'd3045, 32'd3105},
{-32'd6694, 32'd3778, 32'd5802, 32'd3413},
{32'd3354, 32'd3343, -32'd10914, 32'd6738},
{32'd3599, -32'd4385, -32'd893, 32'd17854},
{32'd7986, -32'd4187, 32'd2755, 32'd4981},
{-32'd4842, 32'd4134, 32'd4788, 32'd7830},
{32'd10228, 32'd8340, 32'd360, -32'd16682},
{-32'd5825, -32'd38, -32'd9294, -32'd12439},
{-32'd2292, -32'd2421, -32'd9699, -32'd5860},
{32'd4518, -32'd8094, 32'd7940, -32'd5120},
{-32'd6113, 32'd4593, 32'd14525, -32'd2261},
{-32'd8248, -32'd2566, -32'd8979, -32'd4608},
{-32'd4815, -32'd3558, 32'd9015, 32'd9528},
{-32'd880, -32'd3126, -32'd386, 32'd4847},
{32'd5138, 32'd2135, -32'd10529, -32'd415},
{-32'd9967, -32'd15553, -32'd1458, -32'd789},
{-32'd2768, 32'd1418, -32'd2220, -32'd5722},
{32'd2018, 32'd194, -32'd3521, -32'd2063},
{32'd1005, 32'd269, 32'd5057, 32'd808},
{-32'd10971, -32'd1853, -32'd533, 32'd525},
{32'd5784, -32'd3890, 32'd810, 32'd4416},
{-32'd563, 32'd3868, -32'd3570, 32'd1325},
{32'd2835, 32'd11, -32'd1642, 32'd4820},
{32'd3936, 32'd9107, -32'd185, -32'd204},
{32'd12811, 32'd4081, -32'd638, 32'd6189},
{32'd7875, 32'd9036, 32'd8365, 32'd4044},
{32'd5364, -32'd10699, -32'd8011, -32'd2376},
{-32'd612, -32'd10574, 32'd742, -32'd994},
{-32'd1726, 32'd4707, -32'd2625, 32'd3621},
{-32'd5392, -32'd12984, 32'd1426, -32'd8218},
{-32'd4388, -32'd2741, -32'd6066, 32'd1827},
{-32'd14552, 32'd7748, -32'd7106, -32'd464},
{-32'd5903, 32'd3062, -32'd9782, 32'd848},
{-32'd11134, -32'd1864, -32'd798, -32'd1758},
{-32'd16866, -32'd23032, 32'd1261, -32'd4458},
{-32'd2301, -32'd12281, 32'd12791, 32'd6242},
{32'd1137, -32'd6181, -32'd6249, 32'd3110},
{32'd2944, -32'd4997, 32'd349, 32'd11232},
{32'd4867, 32'd18730, -32'd4082, -32'd10162},
{32'd2750, -32'd12940, -32'd6575, 32'd4317},
{32'd3364, 32'd11395, -32'd8633, 32'd4212},
{32'd1190, -32'd3534, -32'd6696, 32'd6479},
{-32'd496, 32'd331, 32'd1670, 32'd10319},
{32'd8964, -32'd5692, -32'd10917, 32'd6910},
{32'd2065, -32'd5814, -32'd775, 32'd1490},
{32'd1791, -32'd771, -32'd57, -32'd6431},
{-32'd906, 32'd2810, -32'd8042, 32'd209},
{-32'd9813, 32'd10933, 32'd14308, -32'd2797},
{32'd4011, -32'd5364, -32'd1389, 32'd10354},
{32'd5672, -32'd9578, -32'd10741, -32'd2951},
{-32'd4940, -32'd5175, 32'd572, 32'd3109},
{-32'd13510, 32'd7872, 32'd8649, -32'd1558},
{-32'd6233, 32'd4866, -32'd7943, -32'd3054},
{32'd1781, 32'd2985, 32'd10267, -32'd2267},
{32'd10832, 32'd4702, -32'd6999, -32'd663},
{32'd2613, 32'd1172, 32'd15325, 32'd2394},
{32'd12346, -32'd3064, -32'd1510, -32'd4669},
{32'd7538, -32'd3017, 32'd5726, 32'd754},
{32'd5034, -32'd5081, 32'd614, -32'd7330},
{32'd5969, 32'd3144, 32'd1376, -32'd10037},
{-32'd5656, 32'd4204, 32'd2032, -32'd2484},
{-32'd3393, -32'd11161, 32'd11793, 32'd4901},
{-32'd3216, 32'd4594, -32'd1918, -32'd8991},
{-32'd1437, 32'd9993, 32'd11530, -32'd5837},
{32'd5455, 32'd2117, 32'd1934, -32'd881},
{-32'd6347, 32'd6824, 32'd3854, -32'd5116},
{-32'd890, 32'd2933, 32'd4468, 32'd11736},
{-32'd5641, 32'd3439, 32'd5721, 32'd4819},
{-32'd2757, 32'd953, -32'd162, -32'd4633},
{-32'd16837, -32'd2426, -32'd7135, -32'd8057},
{32'd2902, 32'd375, 32'd2160, 32'd2512},
{32'd5169, -32'd1420, -32'd2187, 32'd3181},
{-32'd5534, 32'd702, 32'd12708, 32'd4256},
{-32'd7252, 32'd3073, 32'd4062, 32'd10668},
{-32'd5743, -32'd550, -32'd2779, 32'd375},
{32'd4341, -32'd5085, -32'd1398, 32'd7203},
{32'd1168, -32'd7204, -32'd310, -32'd9408},
{32'd5681, -32'd7571, -32'd525, -32'd9932},
{32'd1957, 32'd2246, -32'd8348, 32'd7377},
{32'd656, 32'd9210, 32'd3204, 32'd5753},
{32'd11132, 32'd20474, -32'd8908, -32'd10041},
{-32'd3113, -32'd7454, 32'd1205, -32'd12014},
{32'd3522, -32'd736, -32'd2728, -32'd426},
{-32'd4244, 32'd9240, 32'd995, -32'd9575},
{-32'd10898, -32'd7502, 32'd4939, 32'd19992},
{32'd762, -32'd417, -32'd6016, -32'd8955},
{-32'd5134, -32'd8197, -32'd4812, 32'd3191},
{32'd933, -32'd1544, 32'd11145, 32'd5338},
{32'd8274, -32'd15461, -32'd10197, -32'd691},
{-32'd15910, -32'd4800, -32'd2801, 32'd4287},
{-32'd2383, 32'd8506, -32'd1442, 32'd306},
{-32'd4129, -32'd14103, -32'd4194, 32'd10335},
{-32'd11400, 32'd6789, 32'd7219, 32'd15026},
{32'd8822, 32'd4095, -32'd1458, 32'd2410},
{32'd8377, 32'd835, 32'd7086, -32'd3926},
{-32'd7868, -32'd11067, -32'd129, 32'd10777},
{-32'd515, 32'd1823, 32'd3975, -32'd3112},
{-32'd5947, 32'd1720, -32'd52, -32'd6074},
{-32'd3930, 32'd11100, -32'd103, -32'd3176},
{-32'd5863, -32'd1731, -32'd3385, -32'd8631},
{-32'd6029, 32'd6318, 32'd5716, -32'd4733},
{-32'd5822, -32'd4309, 32'd5413, -32'd566},
{32'd4173, -32'd1004, 32'd11153, -32'd3839},
{32'd1786, -32'd12597, 32'd12016, -32'd771},
{32'd6138, -32'd9605, -32'd7432, -32'd8064},
{32'd11178, 32'd5681, 32'd2801, 32'd5112},
{-32'd5139, 32'd8147, 32'd390, -32'd4521},
{32'd17334, 32'd2454, -32'd1064, -32'd9473},
{32'd6086, 32'd362, 32'd6897, -32'd662},
{32'd4083, -32'd12538, -32'd5835, 32'd3692},
{-32'd1262, 32'd944, 32'd3633, -32'd4400},
{-32'd7125, -32'd1585, -32'd8053, 32'd3208},
{32'd6444, -32'd1635, 32'd2898, 32'd4363},
{32'd5012, 32'd3818, -32'd2196, -32'd988},
{-32'd7504, -32'd6018, -32'd2048, 32'd3547},
{32'd1303, -32'd5355, -32'd5677, 32'd4547},
{32'd1687, -32'd1643, -32'd2975, 32'd5836},
{-32'd6350, -32'd11192, -32'd5788, 32'd3546},
{32'd6202, -32'd1280, 32'd1988, 32'd5429},
{-32'd9238, -32'd9086, 32'd6586, 32'd11785},
{32'd3730, 32'd8448, 32'd4348, 32'd11754},
{-32'd1986, 32'd566, 32'd7248, 32'd7319},
{-32'd486, 32'd8178, 32'd5667, -32'd13469},
{-32'd618, 32'd8452, 32'd1067, -32'd5465},
{-32'd2436, -32'd3303, -32'd17985, 32'd5263},
{32'd7758, -32'd4064, -32'd7312, -32'd113},
{32'd1926, -32'd62, -32'd10579, -32'd3527},
{-32'd10947, 32'd3358, -32'd9875, 32'd95},
{32'd7816, 32'd15111, -32'd3290, 32'd6935},
{32'd6373, -32'd4634, 32'd2303, 32'd7537},
{32'd12946, 32'd2564, 32'd2723, -32'd1175},
{32'd1565, 32'd6535, -32'd8209, -32'd18663}
},
{{32'd8411, 32'd2731, 32'd3305, -32'd1910},
{-32'd9512, -32'd3513, -32'd7083, -32'd508},
{-32'd2494, -32'd10468, 32'd5082, 32'd2026},
{-32'd1643, 32'd2094, 32'd1634, 32'd3304},
{32'd5738, 32'd558, 32'd12810, 32'd3619},
{-32'd2810, -32'd1874, 32'd4351, -32'd7087},
{32'd1860, 32'd1884, -32'd2364, -32'd2941},
{32'd1719, -32'd5321, -32'd462, 32'd738},
{32'd7524, 32'd2196, 32'd2374, 32'd4778},
{32'd11227, 32'd7657, 32'd1026, 32'd4633},
{32'd2000, -32'd2442, 32'd2924, -32'd3663},
{-32'd4014, -32'd1048, -32'd909, -32'd1015},
{32'd7898, 32'd8329, 32'd3312, 32'd9036},
{32'd4246, -32'd3577, -32'd2432, 32'd1968},
{-32'd2256, -32'd5347, -32'd694, -32'd1335},
{32'd7243, 32'd590, 32'd5483, -32'd11096},
{32'd3698, -32'd432, 32'd8190, -32'd1082},
{32'd9552, -32'd2259, -32'd7297, -32'd3835},
{32'd9482, 32'd2442, 32'd3234, -32'd4631},
{-32'd7355, 32'd2511, 32'd505, 32'd1179},
{-32'd5465, 32'd1518, -32'd9630, 32'd866},
{-32'd6870, -32'd2513, 32'd647, -32'd4946},
{-32'd7696, 32'd2631, 32'd1026, 32'd793},
{-32'd150, 32'd600, -32'd484, -32'd4825},
{-32'd8092, 32'd5701, -32'd1844, 32'd8580},
{-32'd1680, 32'd2947, 32'd13087, -32'd1481},
{32'd478, -32'd6078, 32'd3109, -32'd1008},
{-32'd2996, -32'd4900, -32'd518, 32'd5383},
{-32'd2720, 32'd10749, 32'd2770, 32'd3436},
{-32'd3271, 32'd219, -32'd2698, 32'd3017},
{32'd7875, -32'd5414, 32'd4189, 32'd5982},
{-32'd4695, -32'd4732, -32'd2304, -32'd4987},
{32'd7570, -32'd1028, 32'd7336, 32'd3988},
{32'd3430, -32'd4684, 32'd2952, 32'd199},
{32'd7343, 32'd6414, 32'd4404, 32'd2744},
{32'd2779, 32'd4285, -32'd3036, 32'd3196},
{32'd3055, -32'd2657, 32'd5516, 32'd1443},
{-32'd1341, 32'd860, 32'd3443, 32'd4258},
{32'd4410, 32'd2219, -32'd4766, -32'd3370},
{-32'd348, -32'd7879, -32'd103, -32'd9114},
{-32'd6578, 32'd3659, 32'd7209, -32'd1510},
{32'd3635, -32'd4769, 32'd207, -32'd8161},
{32'd4285, -32'd1058, 32'd8872, -32'd5716},
{-32'd5409, -32'd8281, -32'd5216, -32'd4502},
{32'd9042, -32'd1139, -32'd5976, -32'd2454},
{32'd2888, 32'd5894, -32'd12509, -32'd7107},
{-32'd6602, -32'd1923, -32'd4864, -32'd3746},
{32'd1963, -32'd2788, 32'd2892, -32'd3535},
{-32'd9383, 32'd3969, 32'd4829, 32'd1803},
{-32'd2493, -32'd1363, -32'd14689, -32'd921},
{32'd12077, 32'd606, -32'd561, 32'd2716},
{32'd2886, -32'd4684, -32'd5571, -32'd59},
{-32'd469, 32'd4243, 32'd5035, -32'd3612},
{32'd3631, 32'd6021, -32'd1625, 32'd7123},
{32'd4649, 32'd7448, 32'd3860, -32'd8036},
{32'd2036, -32'd7311, -32'd4662, -32'd1835},
{32'd1322, -32'd8596, 32'd8535, -32'd362},
{32'd3635, 32'd2877, 32'd4107, -32'd10738},
{-32'd5442, -32'd4216, -32'd1517, 32'd1541},
{-32'd5622, -32'd1557, 32'd2006, -32'd931},
{32'd994, -32'd1338, -32'd1175, 32'd8851},
{-32'd6370, 32'd250, 32'd1022, -32'd4259},
{-32'd9011, -32'd4783, -32'd1350, -32'd811},
{-32'd4196, -32'd1127, -32'd2020, -32'd3360},
{32'd2285, 32'd14719, -32'd944, -32'd3362},
{32'd4091, -32'd5233, -32'd4215, 32'd4417},
{-32'd1681, 32'd2483, 32'd3850, -32'd3470},
{-32'd6670, -32'd9855, 32'd1482, 32'd2197},
{-32'd5993, -32'd4838, -32'd12597, 32'd679},
{-32'd5037, -32'd2192, -32'd2263, -32'd3975},
{-32'd638, 32'd775, -32'd9615, -32'd7115},
{32'd133, -32'd4371, -32'd1323, -32'd3418},
{-32'd6111, -32'd7629, -32'd5351, -32'd2625},
{32'd5341, -32'd4436, -32'd4820, -32'd5930},
{-32'd355, 32'd735, 32'd2624, 32'd1728},
{32'd15641, -32'd9867, -32'd8975, -32'd7506},
{-32'd5614, 32'd3206, -32'd2543, -32'd5257},
{32'd322, -32'd940, 32'd2499, -32'd630},
{-32'd2758, 32'd3789, -32'd1580, 32'd1984},
{32'd2651, -32'd3926, 32'd5090, -32'd4887},
{32'd1409, 32'd7061, 32'd2091, -32'd817},
{32'd12667, 32'd3606, -32'd2676, 32'd6074},
{-32'd11168, -32'd475, -32'd2901, -32'd845},
{-32'd1113, -32'd2749, 32'd6027, 32'd2648},
{32'd7644, 32'd2111, -32'd7935, 32'd5253},
{32'd8645, -32'd5981, 32'd3020, -32'd7181},
{-32'd4346, -32'd131, 32'd3664, 32'd2072},
{-32'd9897, 32'd329, -32'd2685, -32'd1324},
{-32'd4116, 32'd7512, 32'd2075, -32'd11},
{-32'd7261, 32'd2633, 32'd4035, -32'd4864},
{32'd3706, 32'd2636, -32'd6510, 32'd2020},
{-32'd8097, -32'd6755, -32'd1953, -32'd6881},
{32'd2897, 32'd7507, 32'd2936, 32'd4808},
{32'd3164, 32'd5090, 32'd6288, 32'd6795},
{32'd4512, -32'd1818, 32'd6973, 32'd1881},
{32'd2400, 32'd228, 32'd10453, -32'd510},
{32'd12182, 32'd3767, 32'd7469, -32'd3087},
{32'd5568, 32'd170, 32'd5585, 32'd8735},
{32'd709, -32'd14651, -32'd5101, -32'd1335},
{32'd6684, 32'd5014, 32'd3686, 32'd1307},
{-32'd4162, 32'd3607, 32'd7320, 32'd1331},
{-32'd5880, 32'd2977, -32'd3141, -32'd4373},
{-32'd7980, -32'd3529, 32'd2197, -32'd5460},
{32'd5572, 32'd13039, -32'd6669, -32'd33},
{32'd1551, -32'd8878, 32'd2618, 32'd6129},
{-32'd1405, 32'd1155, 32'd531, -32'd7723},
{32'd3937, -32'd10037, 32'd3052, 32'd1523},
{32'd3313, 32'd531, -32'd2059, 32'd1327},
{32'd1239, 32'd2091, 32'd3043, 32'd4224},
{32'd3029, 32'd481, 32'd4561, 32'd2503},
{32'd6400, 32'd14841, -32'd780, -32'd1700},
{32'd2000, 32'd4627, 32'd2307, -32'd8943},
{32'd1953, 32'd4247, -32'd2744, 32'd782},
{-32'd2590, 32'd559, -32'd795, 32'd3813},
{-32'd1369, 32'd9027, 32'd6951, 32'd3331},
{-32'd941, 32'd2078, 32'd0, 32'd990},
{32'd934, 32'd13339, 32'd2007, 32'd1687},
{-32'd261, 32'd7268, 32'd503, -32'd4583},
{32'd12746, 32'd5663, -32'd546, 32'd1580},
{32'd15063, 32'd1057, 32'd3388, 32'd7969},
{-32'd4886, -32'd1360, -32'd2247, -32'd1836},
{32'd2116, 32'd3369, 32'd4928, -32'd587},
{32'd6558, -32'd7347, -32'd2700, 32'd5968},
{-32'd8923, -32'd544, 32'd3096, 32'd3396},
{-32'd4445, -32'd2302, 32'd4329, -32'd2710},
{32'd694, 32'd3196, 32'd462, 32'd5959},
{32'd1166, 32'd4672, 32'd4537, -32'd4308},
{-32'd3561, -32'd6036, -32'd7889, 32'd1761},
{-32'd4034, 32'd1200, 32'd4686, -32'd1802},
{32'd4272, 32'd503, -32'd7305, -32'd281},
{-32'd741, 32'd2217, 32'd5395, 32'd1181},
{32'd3158, -32'd4262, -32'd9564, -32'd6194},
{-32'd6384, 32'd2979, -32'd5305, -32'd5296},
{32'd292, -32'd7753, 32'd1755, 32'd5042},
{-32'd7234, -32'd7721, -32'd188, 32'd3732},
{-32'd3059, -32'd2856, -32'd4496, -32'd3178},
{32'd4892, -32'd3875, 32'd1130, -32'd507},
{32'd3879, 32'd1959, -32'd7590, -32'd1980},
{32'd7538, 32'd259, 32'd2095, 32'd2015},
{-32'd11084, -32'd3802, -32'd5287, 32'd508},
{32'd6404, -32'd1488, 32'd6561, 32'd3669},
{32'd10087, -32'd746, 32'd3763, -32'd9421},
{32'd2212, -32'd3610, 32'd4583, 32'd3664},
{-32'd5697, 32'd2597, 32'd2073, -32'd2161},
{32'd6219, 32'd12453, -32'd2975, 32'd5163},
{32'd4563, 32'd959, 32'd5818, 32'd11372},
{-32'd8889, -32'd11931, 32'd5386, -32'd3036},
{32'd10594, 32'd2601, -32'd3116, 32'd2130},
{32'd3337, 32'd3551, -32'd5587, -32'd3376},
{-32'd2949, -32'd8725, 32'd4369, -32'd1447},
{-32'd6863, -32'd5987, -32'd3208, -32'd5998},
{32'd17, -32'd525, -32'd2068, 32'd2194},
{32'd1976, -32'd2130, 32'd4904, -32'd6181},
{32'd3512, -32'd3172, 32'd4969, -32'd6442},
{-32'd7182, -32'd11187, -32'd4224, -32'd5486},
{32'd1262, -32'd883, 32'd2131, 32'd7487},
{32'd1514, -32'd4880, -32'd3780, 32'd4733},
{-32'd7081, -32'd6290, -32'd7446, -32'd1110},
{32'd5479, 32'd3290, 32'd6802, 32'd5984},
{32'd8879, 32'd1745, 32'd8532, -32'd1207},
{-32'd5461, -32'd7732, -32'd5246, 32'd8045},
{32'd4326, -32'd1423, 32'd5117, 32'd2368},
{-32'd4029, 32'd1748, -32'd1769, 32'd1996},
{32'd6701, -32'd11099, -32'd4143, 32'd2412},
{-32'd3248, 32'd4577, -32'd1050, 32'd2955},
{-32'd17345, -32'd3135, -32'd2015, -32'd6067},
{32'd1604, 32'd5775, 32'd10434, 32'd3512},
{32'd2415, 32'd6129, -32'd11651, -32'd3926},
{32'd6148, -32'd936, 32'd1903, 32'd1032},
{-32'd7226, -32'd4423, 32'd1049, -32'd8832},
{-32'd12481, 32'd206, 32'd619, -32'd1862},
{32'd343, -32'd1555, 32'd7454, -32'd3060},
{32'd8392, 32'd1609, 32'd3100, -32'd1305},
{-32'd503, -32'd2662, 32'd1534, 32'd482},
{32'd4134, 32'd997, -32'd6272, 32'd7114},
{32'd2673, -32'd1281, 32'd2135, 32'd4006},
{-32'd982, 32'd1609, 32'd2444, 32'd1847},
{32'd2257, 32'd7649, -32'd4065, -32'd2797},
{-32'd2754, -32'd6100, 32'd2247, 32'd4872},
{32'd1656, -32'd9915, 32'd1957, -32'd1143},
{32'd3096, 32'd5842, -32'd1204, 32'd1498},
{32'd5696, 32'd1223, 32'd3258, -32'd3008},
{32'd1384, 32'd4360, -32'd3066, -32'd6476},
{32'd4158, -32'd4318, 32'd1083, -32'd4670},
{-32'd2638, 32'd10489, 32'd12679, 32'd6334},
{32'd2958, 32'd6431, 32'd8720, 32'd11512},
{-32'd927, 32'd2601, -32'd9646, 32'd6694},
{32'd9782, -32'd241, -32'd8770, -32'd439},
{-32'd2358, -32'd5032, 32'd1537, 32'd12384},
{32'd5674, 32'd6385, -32'd4451, -32'd3676},
{32'd5162, -32'd647, 32'd198, -32'd3669},
{32'd4040, -32'd2827, -32'd1741, -32'd4337},
{32'd453, 32'd4800, 32'd7915, -32'd1167},
{32'd3495, -32'd7664, 32'd5279, 32'd6725},
{32'd7746, -32'd1859, 32'd1302, -32'd3947},
{32'd5750, 32'd5564, -32'd3073, -32'd1471},
{-32'd5453, 32'd2850, 32'd9370, 32'd276},
{32'd8101, -32'd6968, -32'd1630, 32'd7150},
{-32'd519, 32'd4607, -32'd3287, -32'd1954},
{32'd717, 32'd6098, -32'd4081, 32'd6165},
{-32'd12578, -32'd4774, -32'd3313, -32'd3999},
{-32'd1724, -32'd354, 32'd6440, -32'd13167},
{32'd5438, -32'd6464, -32'd6769, 32'd2937},
{32'd687, -32'd8646, -32'd2217, 32'd3688},
{-32'd1760, -32'd333, -32'd3660, -32'd380},
{-32'd3396, 32'd2203, 32'd2387, 32'd234},
{32'd8875, 32'd2338, 32'd2920, 32'd10846},
{-32'd4137, 32'd2040, -32'd1735, -32'd6920},
{32'd4250, 32'd4146, -32'd1006, 32'd1559},
{32'd4641, 32'd617, 32'd3610, -32'd2771},
{32'd9918, -32'd2729, 32'd4894, -32'd7578},
{32'd4649, 32'd12330, -32'd3940, 32'd6486},
{-32'd5381, -32'd4685, -32'd10192, -32'd6845},
{-32'd2080, 32'd3470, 32'd1591, 32'd3750},
{32'd593, -32'd9453, 32'd2120, -32'd3499},
{-32'd4012, 32'd6755, 32'd3387, -32'd1427},
{-32'd6048, -32'd2296, 32'd3013, 32'd4142},
{-32'd2534, 32'd551, -32'd6106, 32'd4075},
{-32'd10439, -32'd2303, 32'd3691, -32'd1862},
{-32'd4885, -32'd9408, -32'd7721, 32'd2471},
{32'd4160, -32'd5006, -32'd5991, 32'd2603},
{32'd3470, 32'd2641, -32'd1201, 32'd5582},
{32'd5848, -32'd1259, 32'd2257, -32'd2343},
{-32'd2363, 32'd1503, -32'd9475, 32'd304},
{-32'd904, 32'd1017, 32'd7156, -32'd901},
{32'd4946, 32'd258, -32'd4735, 32'd4682},
{32'd838, 32'd4943, -32'd2477, 32'd1103},
{-32'd3112, 32'd359, -32'd614, -32'd4561},
{32'd10391, 32'd6024, 32'd904, 32'd1686},
{-32'd2299, -32'd6305, 32'd5777, 32'd3697},
{-32'd6720, -32'd6850, 32'd5355, -32'd5394},
{32'd3220, -32'd1454, 32'd3382, 32'd1961},
{-32'd2377, -32'd5427, 32'd10600, 32'd2706},
{32'd8209, -32'd3409, -32'd2706, 32'd5289},
{32'd3038, -32'd7102, -32'd2416, 32'd5177},
{32'd5376, -32'd5548, -32'd8137, -32'd3557},
{-32'd2804, -32'd1861, 32'd7839, 32'd4141},
{32'd813, -32'd9564, 32'd10037, 32'd4131},
{-32'd7672, 32'd8635, 32'd2785, -32'd13310},
{-32'd4073, -32'd1101, 32'd1461, -32'd1421},
{-32'd7644, -32'd2466, -32'd1944, -32'd4850},
{-32'd5434, -32'd5251, -32'd1233, -32'd1940},
{-32'd11182, 32'd639, 32'd3376, -32'd2082},
{-32'd3239, 32'd3428, 32'd2061, 32'd1962},
{32'd6283, 32'd2074, 32'd6867, 32'd4459},
{32'd10055, -32'd6231, 32'd9905, -32'd4492},
{32'd239, -32'd4821, 32'd1572, 32'd1183},
{-32'd13526, 32'd5441, -32'd5457, -32'd4744},
{32'd6383, 32'd8086, 32'd5496, 32'd255},
{32'd2598, 32'd1438, -32'd1730, 32'd7732},
{32'd1917, 32'd2167, 32'd4358, 32'd8705},
{32'd4646, -32'd5070, 32'd1898, 32'd4863},
{32'd12255, 32'd5569, 32'd391, -32'd1116},
{-32'd4086, 32'd4613, 32'd5123, 32'd7566},
{32'd1133, -32'd3443, -32'd1348, 32'd403},
{32'd6935, 32'd5319, 32'd6016, -32'd1754},
{-32'd4480, 32'd686, 32'd4761, 32'd16},
{32'd11379, -32'd6780, -32'd6583, -32'd593},
{-32'd5128, -32'd8119, 32'd2844, -32'd2537},
{32'd194, 32'd2188, -32'd1800, -32'd4109},
{-32'd7851, 32'd1556, -32'd3827, 32'd6842},
{-32'd5001, 32'd4547, -32'd9279, -32'd3807},
{-32'd2972, 32'd6342, 32'd2643, -32'd2341},
{32'd2637, -32'd3082, 32'd1885, 32'd878},
{32'd2858, -32'd3017, 32'd4494, -32'd1613},
{32'd169, 32'd5699, 32'd1508, 32'd7354},
{32'd3172, 32'd6942, -32'd8007, 32'd405},
{32'd10, -32'd8969, -32'd2829, 32'd2460},
{-32'd13325, 32'd3094, -32'd3731, -32'd256},
{-32'd8238, 32'd9708, 32'd4446, 32'd1611},
{-32'd3888, 32'd3590, -32'd1056, 32'd5732},
{32'd3978, 32'd1831, -32'd630, 32'd4963},
{32'd4602, 32'd3702, -32'd4140, -32'd4147},
{-32'd3887, -32'd1372, -32'd3394, 32'd2093},
{-32'd8325, -32'd2487, -32'd2096, 32'd518},
{-32'd2139, 32'd4008, -32'd2895, -32'd7138},
{32'd12417, 32'd7451, 32'd4974, 32'd3240},
{32'd5433, 32'd8833, 32'd881, 32'd4008},
{-32'd8499, -32'd5579, -32'd3135, -32'd1004},
{-32'd4392, 32'd1978, 32'd4383, -32'd966},
{32'd1416, 32'd5462, -32'd1719, 32'd4088},
{-32'd3631, -32'd1738, -32'd8897, 32'd8551},
{32'd5776, 32'd309, 32'd3852, -32'd3893},
{-32'd1012, -32'd5489, 32'd3069, 32'd4194},
{32'd6381, -32'd759, 32'd5017, 32'd14479},
{-32'd2770, -32'd2190, -32'd126, 32'd3658},
{-32'd1198, 32'd11122, -32'd2569, 32'd3901},
{-32'd3512, -32'd7799, -32'd5700, -32'd1956},
{-32'd371, -32'd5011, -32'd3796, 32'd3936},
{-32'd2993, -32'd10813, 32'd539, -32'd4693},
{32'd1388, 32'd6543, 32'd2580, 32'd10054},
{32'd6282, -32'd43, -32'd4486, 32'd1668},
{32'd134, 32'd6228, 32'd6499, -32'd5949},
{32'd6530, -32'd486, -32'd11184, 32'd2694},
{-32'd377, -32'd5328, -32'd9857, -32'd1900},
{32'd1512, -32'd8849, 32'd1393, -32'd4084},
{32'd8171, 32'd3557, -32'd3538, -32'd1700},
{-32'd3910, 32'd8960, -32'd6314, -32'd2415},
{32'd9077, 32'd1829, 32'd4161, 32'd1656},
{32'd1520, 32'd6923, -32'd3470, -32'd4844}
},
{{-32'd1227, -32'd3311, 32'd10110, 32'd2285},
{-32'd20302, 32'd1434, 32'd3456, -32'd2623},
{32'd5430, 32'd81, 32'd1258, 32'd11521},
{32'd9448, -32'd12882, 32'd12016, 32'd10672},
{32'd2768, 32'd7672, 32'd573, 32'd3926},
{32'd2729, -32'd5099, 32'd941, -32'd5453},
{32'd20097, 32'd8082, 32'd160, -32'd2747},
{32'd877, 32'd2196, -32'd364, 32'd4325},
{-32'd7192, -32'd17740, 32'd7793, 32'd12044},
{32'd7990, 32'd9962, 32'd13068, 32'd2933},
{-32'd3590, -32'd6430, -32'd12641, -32'd6162},
{-32'd8014, -32'd11451, -32'd1869, -32'd5308},
{32'd7335, 32'd8734, 32'd11145, 32'd259},
{32'd288, 32'd4461, -32'd4262, 32'd3268},
{32'd2985, 32'd7126, -32'd1492, 32'd3750},
{-32'd1753, -32'd211, -32'd4477, -32'd6769},
{32'd4163, 32'd9660, 32'd8225, -32'd713},
{32'd357, -32'd3709, 32'd2545, 32'd1070},
{32'd1622, -32'd6462, -32'd9715, 32'd15533},
{32'd749, -32'd8007, 32'd525, 32'd3161},
{32'd9245, 32'd2680, 32'd2660, 32'd3431},
{-32'd9325, -32'd6834, -32'd1988, 32'd4094},
{-32'd10493, -32'd3184, 32'd1540, -32'd2384},
{-32'd3431, -32'd9014, 32'd1848, -32'd4556},
{32'd17805, 32'd4274, -32'd4369, -32'd5132},
{-32'd4538, 32'd11635, 32'd6356, -32'd4399},
{-32'd7820, -32'd7919, -32'd3561, -32'd5967},
{32'd9271, 32'd3529, 32'd5141, -32'd5241},
{-32'd7772, -32'd11931, -32'd1926, -32'd1304},
{-32'd4495, -32'd3248, -32'd6443, 32'd9877},
{-32'd1403, 32'd48, 32'd8895, -32'd2319},
{-32'd3822, -32'd3788, -32'd6554, -32'd4981},
{32'd4692, -32'd3984, -32'd2761, 32'd1383},
{32'd3128, 32'd2993, 32'd1475, -32'd4314},
{32'd1372, 32'd7893, 32'd5500, 32'd3104},
{-32'd1745, -32'd3562, 32'd5704, 32'd6545},
{32'd1798, -32'd6871, -32'd7063, 32'd6628},
{32'd150, 32'd8564, -32'd2729, 32'd6075},
{-32'd12136, -32'd1276, 32'd5313, -32'd649},
{32'd1409, -32'd12099, -32'd6275, 32'd3031},
{-32'd10639, -32'd9000, -32'd10981, -32'd3742},
{32'd5302, -32'd982, -32'd397, 32'd5468},
{-32'd11168, -32'd7606, -32'd10131, -32'd11011},
{32'd5579, 32'd8442, -32'd7010, 32'd3086},
{-32'd231, 32'd6446, 32'd4585, -32'd9526},
{-32'd5329, 32'd2453, -32'd2708, -32'd1631},
{32'd6469, -32'd265, 32'd4865, -32'd2131},
{32'd4655, -32'd12349, 32'd2862, -32'd3456},
{32'd18481, -32'd3443, 32'd8658, -32'd1847},
{-32'd4565, -32'd5367, -32'd6154, -32'd5472},
{-32'd16498, -32'd3155, 32'd10400, -32'd2755},
{32'd203, 32'd5703, -32'd7190, 32'd2727},
{-32'd8528, -32'd11094, -32'd4431, 32'd222},
{-32'd2366, 32'd2366, -32'd2685, 32'd425},
{32'd6086, 32'd1626, -32'd387, -32'd9887},
{-32'd12699, -32'd10198, -32'd6351, 32'd15289},
{32'd7654, 32'd4114, 32'd12261, 32'd5758},
{32'd4314, -32'd4732, -32'd3347, -32'd765},
{-32'd12807, 32'd9114, -32'd11077, -32'd6104},
{-32'd5861, -32'd15690, -32'd1811, -32'd6464},
{-32'd3359, -32'd182, -32'd5559, 32'd7328},
{32'd1338, -32'd411, -32'd6922, 32'd3405},
{-32'd6116, -32'd6037, -32'd490, -32'd8048},
{-32'd17054, 32'd4448, 32'd3669, 32'd8100},
{32'd6207, 32'd13389, -32'd2304, -32'd2047},
{32'd7383, -32'd5396, 32'd11270, 32'd8867},
{-32'd13333, 32'd7671, -32'd3535, -32'd10723},
{-32'd5172, -32'd3200, 32'd4263, 32'd3934},
{-32'd7397, 32'd4912, 32'd1409, 32'd6885},
{32'd1893, 32'd3151, 32'd697, 32'd3432},
{32'd8247, 32'd4522, 32'd1455, -32'd3263},
{-32'd4524, -32'd455, 32'd3718, 32'd1125},
{32'd2826, 32'd8059, -32'd1646, 32'd3203},
{-32'd123, -32'd10383, 32'd3945, -32'd2737},
{32'd4517, -32'd3103, 32'd98, 32'd8508},
{-32'd3369, 32'd8891, 32'd4334, -32'd3868},
{-32'd13480, -32'd9047, -32'd2248, -32'd5030},
{-32'd2612, 32'd2127, -32'd4610, -32'd4969},
{32'd11956, 32'd8930, 32'd9347, 32'd8346},
{-32'd1847, -32'd3056, -32'd2304, 32'd8996},
{-32'd14078, 32'd2878, -32'd3648, 32'd4255},
{32'd3014, 32'd3165, 32'd10306, 32'd7411},
{-32'd10276, -32'd17657, -32'd10934, -32'd1424},
{-32'd6948, 32'd1074, -32'd3277, -32'd1409},
{-32'd9945, -32'd860, -32'd5057, -32'd3774},
{-32'd4568, -32'd11609, 32'd3423, -32'd2242},
{-32'd5594, -32'd3204, 32'd2553, 32'd4412},
{-32'd14863, -32'd5719, -32'd1154, 32'd965},
{-32'd13947, 32'd6746, 32'd6641, 32'd1656},
{-32'd9401, -32'd4657, -32'd2472, -32'd876},
{32'd2437, 32'd9316, 32'd7808, -32'd3081},
{-32'd1219, 32'd1487, -32'd3312, 32'd293},
{32'd15273, 32'd9891, 32'd4781, 32'd8354},
{32'd10991, 32'd11474, 32'd6260, 32'd1472},
{-32'd6138, -32'd775, -32'd7334, -32'd10316},
{-32'd15679, -32'd613, -32'd553, -32'd5527},
{-32'd3136, 32'd8110, 32'd7808, 32'd2919},
{32'd11882, 32'd1747, 32'd3440, 32'd3953},
{-32'd9909, -32'd4070, -32'd1802, 32'd11468},
{32'd7356, 32'd7129, 32'd5652, 32'd4324},
{32'd502, -32'd8421, -32'd11149, -32'd2971},
{-32'd14153, -32'd6618, 32'd4604, -32'd6741},
{-32'd15698, 32'd5364, 32'd8562, 32'd3005},
{-32'd7897, -32'd6766, 32'd4465, -32'd9248},
{-32'd6974, 32'd10941, 32'd6147, -32'd2501},
{-32'd2681, -32'd88, -32'd2314, -32'd120},
{32'd4975, 32'd3764, 32'd4485, -32'd1166},
{32'd3435, 32'd2422, -32'd383, -32'd8753},
{-32'd2834, -32'd384, 32'd5010, -32'd5155},
{-32'd12599, -32'd1072, 32'd6687, 32'd4593},
{-32'd5645, 32'd1001, -32'd1088, 32'd6952},
{-32'd20769, -32'd4761, -32'd1716, 32'd886},
{32'd4565, 32'd16217, 32'd12848, 32'd546},
{32'd18144, 32'd3370, -32'd4015, -32'd6408},
{-32'd7797, -32'd12722, -32'd5246, -32'd4619},
{-32'd3390, -32'd5276, 32'd7787, 32'd9046},
{32'd1546, -32'd240, 32'd10732, -32'd1507},
{-32'd4383, -32'd2473, -32'd2492, -32'd10023},
{32'd6751, 32'd4446, 32'd2770, -32'd9004},
{32'd7305, 32'd5823, 32'd8892, 32'd1025},
{32'd8531, 32'd4545, 32'd8215, 32'd7889},
{-32'd6404, -32'd1797, -32'd222, 32'd15268},
{32'd1831, -32'd2165, 32'd438, -32'd4112},
{32'd442, -32'd113, -32'd3395, -32'd9395},
{-32'd981, -32'd8840, -32'd4713, -32'd2379},
{-32'd10317, 32'd4937, 32'd14315, 32'd7895},
{-32'd1154, -32'd3921, -32'd16318, -32'd8439},
{32'd8104, -32'd8469, 32'd1594, 32'd4763},
{-32'd8121, -32'd7463, -32'd149, 32'd2202},
{-32'd2160, 32'd3153, 32'd236, -32'd1694},
{-32'd4110, 32'd4770, 32'd2735, 32'd10806},
{-32'd7115, 32'd10116, -32'd7598, -32'd5485},
{32'd3383, -32'd1678, -32'd6501, -32'd2803},
{32'd12249, 32'd342, -32'd1484, 32'd889},
{32'd10598, -32'd436, 32'd3436, 32'd9337},
{32'd8162, -32'd1292, -32'd4282, -32'd589},
{32'd4611, -32'd3424, 32'd3427, 32'd8917},
{-32'd15711, -32'd10158, 32'd7779, 32'd8467},
{-32'd3775, 32'd4903, -32'd6220, -32'd4108},
{-32'd5120, -32'd4384, 32'd1793, -32'd13107},
{-32'd8418, -32'd4675, 32'd1019, -32'd86},
{32'd1595, 32'd457, -32'd3210, -32'd1945},
{32'd5402, -32'd1061, -32'd2567, 32'd9125},
{32'd12464, 32'd599, -32'd1443, 32'd717},
{32'd1110, -32'd6626, 32'd5198, 32'd9738},
{32'd8794, 32'd2784, 32'd4261, 32'd1430},
{32'd3036, -32'd6014, -32'd7810, -32'd1829},
{32'd2627, -32'd12850, -32'd6463, 32'd6730},
{32'd9123, -32'd2347, 32'd12500, 32'd9054},
{32'd1115, -32'd8397, 32'd5205, 32'd999},
{32'd10380, 32'd3768, -32'd4576, -32'd401},
{-32'd1915, 32'd2582, 32'd2090, 32'd1983},
{-32'd7920, -32'd5336, -32'd687, -32'd7296},
{-32'd3465, 32'd7592, -32'd3474, -32'd207},
{-32'd7432, -32'd7181, -32'd1494, 32'd4304},
{32'd7031, 32'd9079, 32'd6427, -32'd136},
{32'd7575, -32'd2246, -32'd1092, 32'd12117},
{32'd3021, 32'd4423, 32'd7306, -32'd8144},
{-32'd10479, -32'd3911, 32'd651, -32'd3286},
{-32'd8935, 32'd14806, 32'd1961, 32'd6924},
{32'd3749, 32'd13541, 32'd5613, -32'd4198},
{32'd517, -32'd231, 32'd5550, 32'd10457},
{-32'd6653, -32'd2525, -32'd6886, -32'd3613},
{32'd12680, 32'd5440, 32'd2452, 32'd5531},
{32'd6640, -32'd6775, -32'd586, 32'd4436},
{-32'd3122, 32'd726, -32'd3284, 32'd30},
{32'd755, 32'd8295, 32'd5061, -32'd4566},
{-32'd6807, -32'd5872, -32'd441, 32'd3376},
{32'd7965, 32'd13472, -32'd7365, -32'd2379},
{32'd8467, -32'd6679, -32'd7265, -32'd5698},
{-32'd3694, -32'd11247, 32'd92, -32'd3207},
{32'd2115, -32'd8955, -32'd5708, -32'd1196},
{-32'd1077, 32'd11608, 32'd5765, -32'd1097},
{32'd12653, -32'd4645, -32'd5864, -32'd9047},
{32'd2266, 32'd5363, 32'd9846, 32'd6201},
{-32'd9020, 32'd10989, 32'd454, 32'd9045},
{32'd6226, 32'd3929, 32'd2106, -32'd4438},
{32'd10306, -32'd7795, 32'd4376, 32'd1356},
{32'd5800, 32'd6648, 32'd15752, 32'd10904},
{32'd3977, -32'd248, -32'd7558, -32'd3689},
{32'd3463, -32'd1141, 32'd7726, -32'd13223},
{-32'd2743, 32'd1414, -32'd10559, 32'd6014},
{-32'd2222, -32'd12361, -32'd16190, -32'd14017},
{32'd7743, -32'd5152, -32'd5549, 32'd9138},
{-32'd3856, 32'd8040, 32'd3694, -32'd6120},
{32'd3877, -32'd1487, -32'd8395, -32'd2084},
{-32'd1029, -32'd1842, 32'd5060, -32'd367},
{32'd5126, -32'd5133, 32'd5904, 32'd1978},
{-32'd4148, -32'd3929, -32'd193, -32'd3855},
{32'd722, 32'd11631, -32'd10975, -32'd7356},
{32'd6771, 32'd8308, -32'd5080, -32'd2652},
{32'd6028, 32'd8836, -32'd1418, -32'd10644},
{-32'd8191, -32'd12734, -32'd7914, -32'd4253},
{32'd9291, 32'd7331, 32'd1463, 32'd15018},
{-32'd1114, -32'd4087, 32'd4897, 32'd5010},
{-32'd11601, -32'd12617, -32'd7559, -32'd1792},
{-32'd13998, 32'd11950, -32'd5768, -32'd6661},
{-32'd507, -32'd373, 32'd2567, -32'd4883},
{32'd2436, -32'd2496, 32'd2112, 32'd2347},
{32'd3445, -32'd2144, -32'd1398, -32'd9218},
{-32'd3678, -32'd3443, -32'd7073, -32'd2282},
{-32'd3750, -32'd6521, -32'd10967, -32'd8613},
{-32'd4676, -32'd9119, 32'd4656, 32'd4623},
{-32'd3915, 32'd5031, 32'd6207, -32'd11824},
{-32'd7656, -32'd1748, -32'd6093, 32'd8046},
{-32'd5695, 32'd4208, -32'd2323, -32'd2387},
{32'd4097, -32'd691, -32'd7051, 32'd8845},
{-32'd12065, -32'd18999, 32'd6674, -32'd5217},
{32'd2536, 32'd4174, -32'd640, 32'd10916},
{-32'd7300, -32'd8501, -32'd4516, -32'd808},
{-32'd1056, 32'd2059, 32'd6089, -32'd994},
{32'd2338, 32'd10360, 32'd7418, -32'd8986},
{-32'd6333, -32'd2146, 32'd1050, 32'd1087},
{-32'd15062, -32'd3704, 32'd3113, 32'd3044},
{32'd1707, 32'd4374, -32'd5154, -32'd8669},
{-32'd4770, -32'd2054, -32'd4893, -32'd1017},
{-32'd5275, 32'd570, 32'd2074, 32'd5559},
{32'd2912, -32'd11021, 32'd2109, -32'd6341},
{-32'd226, 32'd5129, -32'd667, -32'd6228},
{32'd5598, -32'd1760, -32'd1907, -32'd1538},
{32'd2262, 32'd1755, 32'd8461, -32'd2016},
{32'd2950, 32'd890, 32'd1674, -32'd1436},
{32'd5141, 32'd8948, 32'd5272, 32'd6978},
{32'd12359, 32'd2438, -32'd7944, 32'd6840},
{-32'd6630, -32'd7635, -32'd2803, 32'd7069},
{-32'd16049, 32'd2725, 32'd12800, 32'd3083},
{-32'd8915, 32'd409, -32'd3142, 32'd7012},
{-32'd16318, -32'd11331, -32'd6389, 32'd1618},
{-32'd9494, -32'd3433, -32'd461, 32'd3642},
{32'd3772, -32'd448, 32'd2962, 32'd2506},
{-32'd4462, -32'd2262, -32'd1099, -32'd6699},
{32'd1602, 32'd2934, -32'd206, 32'd202},
{-32'd5058, -32'd1605, 32'd3275, -32'd1028},
{-32'd1387, 32'd3752, 32'd3171, -32'd3481},
{32'd13769, 32'd6004, -32'd14809, -32'd362},
{-32'd194, -32'd3698, -32'd6466, 32'd9023},
{32'd1586, 32'd7402, 32'd2816, 32'd6812},
{32'd3144, 32'd4529, 32'd6822, -32'd12599},
{32'd1874, -32'd5650, -32'd9910, -32'd7487},
{-32'd14160, -32'd9558, -32'd8982, 32'd5867},
{32'd1611, -32'd9098, 32'd399, 32'd3271},
{-32'd10960, -32'd2551, 32'd10442, 32'd683},
{-32'd885, 32'd1846, -32'd2689, -32'd4659},
{32'd4608, 32'd2860, 32'd513, -32'd3978},
{32'd4936, 32'd8538, 32'd4080, 32'd4943},
{-32'd2318, 32'd3250, -32'd8044, -32'd3384},
{32'd6332, 32'd587, -32'd3297, -32'd5394},
{-32'd12394, -32'd6908, 32'd58, -32'd3252},
{32'd10950, 32'd2721, -32'd5272, -32'd9280},
{32'd1411, -32'd830, 32'd5951, -32'd6913},
{-32'd10895, -32'd1367, -32'd7932, -32'd3216},
{32'd9981, 32'd3757, 32'd99, 32'd3156},
{32'd10796, 32'd3952, -32'd5206, -32'd7751},
{32'd14929, 32'd4794, 32'd1918, -32'd753},
{-32'd3615, 32'd1257, -32'd6137, -32'd4382},
{32'd7806, 32'd112, 32'd2625, 32'd2866},
{-32'd3147, -32'd6630, -32'd1852, -32'd1370},
{32'd3452, 32'd14411, 32'd13838, 32'd3325},
{32'd6302, -32'd2686, 32'd2909, -32'd14000},
{-32'd15892, -32'd490, -32'd4939, -32'd4765},
{32'd11392, 32'd3036, 32'd8203, 32'd10361},
{32'd2403, 32'd8384, -32'd3061, 32'd1736},
{-32'd2852, -32'd2750, -32'd7062, 32'd2415},
{-32'd602, 32'd3067, -32'd1403, 32'd8789},
{32'd2198, -32'd4722, 32'd9791, 32'd405},
{-32'd5480, -32'd7976, -32'd1775, -32'd2048},
{32'd14100, -32'd1662, 32'd1672, -32'd1201},
{-32'd8605, -32'd4990, 32'd5623, 32'd7090},
{-32'd3262, 32'd2701, -32'd7006, 32'd1908},
{32'd4526, -32'd11744, -32'd4099, 32'd2036},
{32'd13967, -32'd7974, 32'd1421, -32'd3059},
{-32'd3297, -32'd8165, -32'd2231, 32'd7871},
{-32'd17395, 32'd508, -32'd3160, 32'd3782},
{-32'd5713, 32'd3702, -32'd5971, 32'd3354},
{32'd1990, -32'd2109, 32'd1240, -32'd9077},
{-32'd4654, -32'd8195, -32'd10855, -32'd1364},
{32'd5788, 32'd7483, 32'd8797, 32'd6082},
{32'd7082, -32'd429, -32'd3595, -32'd8163},
{-32'd8065, -32'd13446, -32'd12396, 32'd1363},
{-32'd14248, -32'd9169, -32'd6272, -32'd2688},
{32'd1576, -32'd500, 32'd71, 32'd5907},
{32'd11796, 32'd11851, -32'd6959, -32'd4915},
{32'd8171, 32'd1144, 32'd3992, -32'd3371},
{32'd1355, -32'd9070, 32'd3020, 32'd6666},
{-32'd9144, -32'd11000, 32'd395, -32'd6838},
{32'd7505, -32'd2517, -32'd6360, -32'd12019},
{-32'd108, -32'd4284, 32'd2523, 32'd2359},
{-32'd9750, -32'd4911, -32'd11682, -32'd2199},
{32'd818, 32'd5553, 32'd1663, -32'd4791},
{-32'd10677, -32'd2471, -32'd5316, 32'd1911},
{32'd1121, 32'd5477, 32'd9277, 32'd10451},
{32'd8745, 32'd2019, -32'd1370, 32'd5265},
{-32'd11530, 32'd11267, -32'd2670, -32'd2018},
{-32'd5179, 32'd702, -32'd617, 32'd3462},
{32'd8032, 32'd7113, -32'd2616, -32'd10521},
{32'd6493, 32'd3736, -32'd10643, 32'd547},
{-32'd10628, -32'd11341, -32'd2475, -32'd5517},
{-32'd2728, 32'd871, 32'd880, 32'd4817},
{32'd1884, -32'd15782, -32'd864, -32'd6116},
{32'd119, -32'd694, -32'd623, 32'd3273}
},
{{32'd11814, 32'd1191, -32'd2696, 32'd7022},
{32'd547, -32'd2230, 32'd1367, 32'd833},
{32'd3001, 32'd12998, 32'd3324, 32'd5325},
{-32'd1394, -32'd6754, -32'd2474, -32'd11822},
{-32'd1982, 32'd3542, -32'd974, -32'd9668},
{32'd16146, -32'd1868, 32'd4648, 32'd8252},
{-32'd4970, -32'd10150, -32'd5052, 32'd2243},
{-32'd8847, 32'd2596, -32'd1836, -32'd3172},
{32'd430, 32'd10181, -32'd3344, -32'd4956},
{32'd400, 32'd1036, 32'd1121, -32'd3907},
{32'd5343, 32'd2086, -32'd5538, 32'd2107},
{-32'd182, 32'd5521, 32'd5040, 32'd1078},
{32'd9671, 32'd5940, -32'd3741, 32'd10833},
{32'd415, -32'd10657, 32'd8919, -32'd10870},
{32'd12136, -32'd9955, -32'd8494, -32'd4809},
{32'd6291, 32'd7565, -32'd2201, 32'd9012},
{-32'd13940, 32'd1443, -32'd308, -32'd723},
{-32'd6914, -32'd7357, -32'd3700, 32'd1898},
{32'd2999, -32'd4551, 32'd14751, -32'd10283},
{32'd8987, -32'd113, 32'd3656, 32'd715},
{-32'd17777, 32'd1449, 32'd7611, -32'd11422},
{-32'd3832, -32'd9147, -32'd1206, 32'd10178},
{32'd1980, 32'd4090, 32'd11200, -32'd1843},
{-32'd3620, -32'd3059, 32'd6250, -32'd3169},
{-32'd1531, -32'd7202, 32'd19800, 32'd1677},
{-32'd3400, -32'd2601, -32'd1962, -32'd1859},
{32'd8057, 32'd1917, 32'd2653, 32'd10517},
{32'd2441, 32'd18473, 32'd4256, 32'd7701},
{-32'd8230, 32'd5923, 32'd6853, -32'd4439},
{32'd559, -32'd23284, -32'd2908, 32'd6348},
{-32'd636, 32'd8308, -32'd991, 32'd403},
{32'd8944, -32'd12303, 32'd12408, -32'd8284},
{-32'd12458, 32'd6884, -32'd3144, 32'd2518},
{32'd1054, -32'd1692, -32'd3079, 32'd14419},
{32'd4339, 32'd1168, -32'd2679, -32'd895},
{32'd11323, -32'd675, 32'd1573, -32'd10325},
{-32'd1369, 32'd711, 32'd5611, -32'd281},
{-32'd2640, -32'd10673, 32'd12361, -32'd8512},
{-32'd10001, 32'd192, -32'd3920, 32'd5973},
{32'd5670, -32'd3703, 32'd2726, 32'd11653},
{-32'd10495, -32'd3263, -32'd9795, -32'd5263},
{32'd9701, -32'd10118, -32'd3763, 32'd8334},
{-32'd2806, 32'd415, 32'd15170, 32'd3949},
{32'd12057, -32'd14098, 32'd4459, 32'd3759},
{-32'd2727, 32'd4549, -32'd3469, -32'd2087},
{-32'd368, -32'd6820, 32'd1954, 32'd15312},
{32'd9182, -32'd5910, 32'd6020, -32'd2736},
{-32'd4565, -32'd10320, 32'd2219, -32'd587},
{32'd10895, 32'd14953, -32'd7099, -32'd4524},
{32'd9818, 32'd3377, -32'd8211, -32'd2487},
{-32'd9340, 32'd14419, 32'd14037, 32'd2403},
{32'd9622, -32'd1229, -32'd4342, 32'd6521},
{-32'd5378, 32'd6131, -32'd6133, -32'd6693},
{32'd1587, 32'd341, -32'd1606, -32'd6322},
{-32'd13120, -32'd3173, -32'd5210, -32'd3907},
{32'd3568, 32'd1919, -32'd5306, 32'd3827},
{-32'd7857, -32'd193, -32'd6499, -32'd1336},
{32'd1238, 32'd8662, -32'd1313, 32'd8008},
{-32'd587, 32'd7490, -32'd603, 32'd2308},
{-32'd5266, -32'd5114, 32'd4142, -32'd4209},
{-32'd7383, 32'd2596, 32'd4826, -32'd19311},
{32'd673, -32'd2606, 32'd4728, -32'd1083},
{32'd564, -32'd6190, 32'd3878, -32'd514},
{32'd11964, 32'd4083, -32'd11803, -32'd9727},
{-32'd3749, -32'd489, -32'd12237, 32'd4182},
{32'd2952, -32'd1314, 32'd3694, 32'd1989},
{-32'd5949, -32'd5081, -32'd2025, -32'd7205},
{-32'd3139, 32'd717, -32'd2650, 32'd5396},
{-32'd488, 32'd5011, -32'd510, 32'd2889},
{32'd7527, -32'd8427, -32'd560, 32'd4322},
{-32'd8518, 32'd10047, -32'd6401, 32'd1381},
{32'd18499, -32'd3406, 32'd16188, 32'd10142},
{32'd3669, -32'd11708, -32'd5665, 32'd15637},
{-32'd9266, 32'd49, -32'd3708, -32'd4380},
{-32'd7576, -32'd1237, -32'd10089, -32'd3428},
{32'd5590, 32'd2304, -32'd1645, 32'd6692},
{-32'd14666, -32'd8080, 32'd2728, 32'd2620},
{-32'd7904, -32'd12668, -32'd7491, 32'd4690},
{32'd8953, 32'd2907, 32'd4213, -32'd4128},
{-32'd3341, 32'd7603, -32'd3726, 32'd6866},
{-32'd4691, 32'd11558, -32'd2266, -32'd4442},
{32'd5767, -32'd6023, -32'd7902, -32'd5119},
{-32'd10302, 32'd8064, 32'd6658, 32'd9700},
{-32'd5472, 32'd6921, -32'd5791, 32'd9365},
{-32'd3382, -32'd5511, 32'd11056, -32'd260},
{32'd10536, -32'd1022, 32'd6648, -32'd2997},
{-32'd563, -32'd4424, -32'd2830, 32'd3973},
{-32'd16076, -32'd357, 32'd2235, -32'd1302},
{-32'd12013, 32'd11398, -32'd7424, 32'd1808},
{-32'd9098, 32'd1836, -32'd5452, -32'd8055},
{32'd4349, 32'd200, 32'd10666, -32'd1588},
{-32'd3194, -32'd13880, -32'd4266, -32'd9112},
{-32'd1774, 32'd3911, -32'd1943, -32'd1208},
{-32'd4220, -32'd1965, -32'd9577, -32'd13129},
{-32'd327, 32'd301, 32'd5808, -32'd5255},
{-32'd9847, 32'd5274, -32'd7382, -32'd4585},
{-32'd7769, -32'd937, 32'd5468, -32'd11169},
{32'd1656, -32'd574, 32'd6419, 32'd1060},
{-32'd2060, 32'd3266, 32'd2051, -32'd4909},
{-32'd2291, 32'd9808, 32'd2024, 32'd2966},
{32'd6330, 32'd1198, 32'd1261, -32'd12121},
{32'd4838, -32'd5908, 32'd4407, 32'd9359},
{32'd9235, 32'd1198, 32'd3205, -32'd7605},
{32'd471, -32'd2824, 32'd1699, 32'd4781},
{32'd5232, 32'd8729, 32'd1250, 32'd5230},
{32'd2012, 32'd12438, -32'd3395, -32'd15002},
{32'd9060, -32'd6380, -32'd4052, -32'd5462},
{-32'd1581, -32'd2972, 32'd7723, 32'd236},
{-32'd12961, -32'd8169, 32'd12917, -32'd3385},
{-32'd5044, -32'd2519, 32'd14449, 32'd5618},
{-32'd14220, 32'd15270, -32'd9624, 32'd7811},
{-32'd8944, 32'd7241, 32'd9779, 32'd8506},
{-32'd1949, -32'd12877, -32'd3527, -32'd2746},
{32'd7179, 32'd3513, 32'd5700, 32'd1550},
{32'd9300, -32'd215, -32'd4803, 32'd2533},
{32'd6754, -32'd4759, 32'd850, -32'd3661},
{32'd2179, 32'd3514, -32'd1607, -32'd1094},
{32'd12280, 32'd2904, 32'd1855, 32'd16488},
{-32'd7498, -32'd8981, 32'd4182, -32'd11261},
{32'd11201, -32'd2747, -32'd5529, -32'd1722},
{32'd10089, -32'd3807, 32'd6448, -32'd1248},
{32'd132, 32'd9683, 32'd2166, -32'd6736},
{-32'd2998, 32'd2889, -32'd18933, 32'd7904},
{32'd3697, -32'd8889, 32'd9258, -32'd7730},
{32'd2055, -32'd2430, 32'd3005, -32'd16992},
{-32'd9925, 32'd6997, -32'd9011, -32'd3154},
{32'd7408, -32'd1598, 32'd4837, -32'd1442},
{-32'd17013, 32'd16420, -32'd8481, 32'd1737},
{32'd11967, 32'd6315, 32'd795, 32'd11150},
{-32'd11005, 32'd9344, 32'd5461, 32'd1363},
{-32'd547, -32'd8188, 32'd2879, 32'd5430},
{32'd2925, 32'd2833, 32'd10079, 32'd7482},
{-32'd9590, -32'd5644, -32'd1613, 32'd610},
{-32'd2515, 32'd5112, -32'd10592, -32'd8462},
{-32'd2334, 32'd12735, 32'd22439, 32'd2850},
{32'd6710, 32'd6120, 32'd3897, 32'd13833},
{32'd777, 32'd5288, 32'd140, 32'd12072},
{-32'd407, -32'd4108, 32'd6783, -32'd76},
{32'd18823, 32'd7739, 32'd15662, 32'd9477},
{32'd10104, 32'd56, 32'd434, -32'd4566},
{-32'd1056, 32'd10116, 32'd9104, 32'd602},
{-32'd10505, -32'd2679, -32'd544, 32'd6225},
{-32'd2640, -32'd11951, -32'd8490, -32'd2700},
{32'd18013, 32'd6925, 32'd9207, -32'd10776},
{-32'd37, -32'd3307, 32'd5148, -32'd11648},
{32'd6635, 32'd7804, -32'd5421, 32'd3845},
{-32'd5284, -32'd1500, 32'd815, 32'd1291},
{-32'd10480, -32'd3785, 32'd10542, 32'd9162},
{32'd1000, -32'd12838, 32'd489, -32'd10624},
{-32'd4639, -32'd11162, -32'd1506, 32'd5779},
{32'd8447, 32'd5475, -32'd6539, 32'd7303},
{-32'd2802, 32'd4053, -32'd19493, -32'd4497},
{32'd6527, 32'd3096, -32'd3130, 32'd6513},
{-32'd591, -32'd3955, -32'd8614, 32'd9423},
{-32'd12602, -32'd9068, 32'd2288, 32'd7190},
{-32'd10388, 32'd9227, 32'd1072, -32'd12796},
{-32'd3431, -32'd3350, 32'd6978, -32'd1115},
{-32'd3003, -32'd4375, 32'd1901, -32'd2590},
{-32'd13011, -32'd4375, -32'd6571, -32'd4113},
{32'd7185, 32'd159, 32'd14533, 32'd274},
{32'd4767, 32'd1567, 32'd4379, 32'd363},
{-32'd5780, 32'd2988, 32'd3193, -32'd5341},
{-32'd9114, -32'd3931, 32'd11115, -32'd6162},
{32'd4635, 32'd8563, -32'd4283, -32'd5708},
{32'd3245, -32'd13519, 32'd10258, -32'd3733},
{-32'd1671, -32'd14471, -32'd4776, 32'd5738},
{32'd1862, 32'd52, -32'd9369, -32'd2751},
{-32'd1597, 32'd2070, 32'd7594, 32'd6448},
{32'd940, 32'd2225, 32'd4627, 32'd8997},
{32'd3966, 32'd1243, 32'd1627, 32'd3405},
{32'd9888, -32'd16434, -32'd453, -32'd4384},
{32'd340, -32'd4782, -32'd4221, 32'd233},
{-32'd3040, 32'd1326, -32'd460, 32'd10092},
{32'd5983, -32'd1864, -32'd8011, -32'd15360},
{32'd15683, -32'd1935, 32'd3547, -32'd15532},
{-32'd6463, 32'd1467, 32'd4085, -32'd2158},
{-32'd4207, 32'd3765, -32'd744, 32'd6069},
{-32'd4295, -32'd119, -32'd1548, -32'd5717},
{-32'd7297, -32'd3361, 32'd14204, -32'd10465},
{32'd2550, 32'd341, -32'd9586, 32'd4209},
{-32'd5509, -32'd8146, 32'd7882, -32'd5498},
{32'd4298, 32'd1028, -32'd9127, 32'd9174},
{-32'd3826, -32'd1439, -32'd4044, 32'd2009},
{32'd6094, 32'd1870, 32'd877, 32'd5699},
{32'd6434, 32'd10409, -32'd10241, -32'd584},
{-32'd4719, 32'd2809, -32'd3908, -32'd5076},
{32'd4237, 32'd864, 32'd10278, -32'd3577},
{-32'd1934, 32'd5056, -32'd2883, 32'd2222},
{-32'd4195, 32'd8070, 32'd2244, -32'd2241},
{32'd6355, 32'd9980, 32'd11123, -32'd4602},
{32'd2418, 32'd9, 32'd1043, 32'd1540},
{32'd14441, -32'd18496, 32'd15447, 32'd8233},
{-32'd4652, -32'd1645, -32'd563, -32'd2111},
{-32'd3320, 32'd2219, 32'd5430, -32'd9593},
{32'd8861, 32'd14189, -32'd15020, 32'd10627},
{32'd8460, 32'd15456, 32'd2687, 32'd4515},
{-32'd577, 32'd3977, 32'd1174, -32'd7430},
{-32'd8800, -32'd1667, 32'd3331, 32'd10416},
{-32'd3297, 32'd7032, -32'd2999, -32'd10573},
{-32'd3718, -32'd1975, 32'd10990, 32'd3910},
{-32'd2167, -32'd1089, -32'd1866, -32'd799},
{32'd2397, 32'd5664, -32'd5214, 32'd4996},
{-32'd2123, 32'd14676, -32'd11129, 32'd3656},
{-32'd10700, -32'd1282, -32'd4015, -32'd1180},
{32'd1318, 32'd2051, 32'd5408, -32'd4045},
{-32'd5960, -32'd9528, -32'd8102, -32'd10081},
{-32'd2523, 32'd9318, -32'd6746, -32'd11162},
{32'd9368, 32'd5519, -32'd5109, -32'd3037},
{-32'd2659, 32'd13986, -32'd3939, -32'd2457},
{32'd3189, 32'd5344, 32'd4112, 32'd3511},
{-32'd5582, 32'd9890, -32'd8627, 32'd5381},
{-32'd1153, -32'd768, -32'd15135, 32'd1499},
{32'd9668, 32'd535, 32'd8270, 32'd2427},
{32'd3963, 32'd2705, -32'd9844, -32'd5614},
{32'd4873, 32'd7106, 32'd8581, 32'd3733},
{32'd3943, 32'd6044, -32'd12432, -32'd8334},
{32'd2640, -32'd3031, -32'd9262, -32'd413},
{-32'd5967, -32'd10422, -32'd7086, 32'd11108},
{32'd518, -32'd9977, -32'd720, -32'd99},
{32'd4205, 32'd5601, 32'd1375, -32'd2563},
{32'd4995, -32'd1688, -32'd2743, 32'd3004},
{32'd3200, -32'd6048, 32'd22384, 32'd528},
{32'd3701, 32'd17760, 32'd1386, -32'd2873},
{32'd2894, -32'd4730, 32'd1460, 32'd3619},
{32'd12465, 32'd532, 32'd3288, -32'd1386},
{32'd1786, -32'd4107, 32'd1428, -32'd8173},
{32'd4229, -32'd1735, -32'd3037, 32'd635},
{-32'd8240, 32'd2992, 32'd6224, -32'd819},
{32'd5318, 32'd4909, 32'd10747, -32'd8400},
{32'd2018, -32'd2263, 32'd6547, 32'd14762},
{32'd89, 32'd2624, 32'd2194, 32'd8932},
{32'd2040, 32'd10913, -32'd1078, -32'd1453},
{32'd7088, 32'd5546, -32'd10285, -32'd2096},
{32'd4065, 32'd16172, 32'd11076, 32'd7692},
{32'd6047, -32'd7403, -32'd9322, 32'd10284},
{-32'd1767, 32'd1216, 32'd1626, 32'd6153},
{32'd1777, -32'd10922, -32'd1989, -32'd1544},
{32'd14238, 32'd4772, -32'd2383, -32'd3039},
{32'd213, 32'd2766, 32'd14479, 32'd13403},
{32'd3841, -32'd2299, 32'd9698, 32'd5824},
{-32'd5836, -32'd11242, -32'd3009, -32'd8802},
{32'd2217, 32'd12641, -32'd1584, 32'd2644},
{32'd5110, 32'd4344, -32'd1129, -32'd225},
{32'd1095, -32'd4131, 32'd2457, -32'd13684},
{-32'd3822, 32'd8996, -32'd556, -32'd3618},
{-32'd4384, 32'd1728, -32'd3719, -32'd6210},
{32'd8804, 32'd2114, -32'd288, 32'd9156},
{32'd2229, -32'd8674, 32'd7624, 32'd1855},
{-32'd5629, 32'd5906, -32'd4633, -32'd9317},
{-32'd2231, -32'd8042, -32'd5921, 32'd3331},
{32'd6242, 32'd495, -32'd11300, -32'd5146},
{32'd782, -32'd5276, -32'd550, -32'd904},
{32'd884, 32'd2300, -32'd117, 32'd6315},
{32'd16305, -32'd2790, -32'd10305, -32'd4319},
{32'd2631, 32'd3572, -32'd2294, -32'd1266},
{-32'd689, 32'd6323, 32'd4465, -32'd9766},
{-32'd6672, 32'd1896, -32'd10342, -32'd12682},
{32'd6473, -32'd864, 32'd6288, -32'd1640},
{-32'd2150, -32'd15235, -32'd5965, 32'd5936},
{32'd1275, -32'd5454, 32'd10785, 32'd6383},
{-32'd3301, -32'd4527, -32'd8543, -32'd7884},
{-32'd5076, -32'd13838, 32'd3601, -32'd2385},
{32'd7536, -32'd1978, -32'd3290, -32'd2013},
{32'd5201, 32'd9436, -32'd3639, 32'd14936},
{-32'd7395, 32'd10287, 32'd1790, 32'd3052},
{-32'd5661, -32'd7808, 32'd3636, -32'd1271},
{32'd12236, -32'd13639, 32'd8082, -32'd7486},
{32'd6022, -32'd11571, 32'd13012, 32'd2076},
{-32'd6068, -32'd10818, 32'd2928, -32'd2195},
{-32'd10173, -32'd2401, -32'd7620, 32'd1580},
{-32'd4538, -32'd5565, 32'd2130, 32'd8695},
{32'd422, 32'd4309, 32'd7448, -32'd7568},
{-32'd12038, 32'd19610, -32'd6720, -32'd311},
{32'd7906, -32'd6729, -32'd1128, 32'd4159},
{32'd8054, -32'd15030, -32'd153, -32'd5112},
{-32'd1414, 32'd5104, -32'd3660, 32'd14545},
{32'd368, 32'd2882, 32'd9057, -32'd3449},
{-32'd5800, -32'd9357, -32'd9851, -32'd1828},
{32'd996, 32'd3186, 32'd3028, 32'd9775},
{32'd7535, -32'd9634, 32'd2241, 32'd7190},
{32'd5550, 32'd7813, 32'd12218, -32'd8023},
{32'd8268, 32'd13076, 32'd2660, -32'd829},
{-32'd16854, 32'd11224, -32'd840, 32'd88},
{32'd1469, -32'd554, -32'd5899, -32'd1598},
{-32'd17816, 32'd3898, 32'd13636, -32'd1216},
{32'd707, -32'd8886, -32'd6908, -32'd3310},
{-32'd3530, 32'd6407, -32'd9133, -32'd1395},
{32'd14596, -32'd1112, -32'd1399, -32'd4071},
{32'd9945, -32'd11309, 32'd9381, -32'd5664},
{32'd2953, 32'd3412, 32'd1494, 32'd8313},
{32'd3235, 32'd1041, 32'd4097, -32'd8710},
{32'd3174, 32'd7945, 32'd18260, -32'd427},
{-32'd4212, 32'd467, -32'd8622, -32'd10314},
{-32'd110, -32'd12958, -32'd859, 32'd9773},
{32'd12613, -32'd1950, 32'd6670, 32'd2132},
{32'd2882, 32'd2109, -32'd2869, 32'd17362},
{32'd7899, 32'd9435, -32'd2768, -32'd11453},
{32'd62, -32'd298, -32'd5825, -32'd1206},
{-32'd3035, 32'd7181, 32'd175, 32'd1162},
{32'd478, -32'd7448, 32'd1374, 32'd8839}
},
{{32'd12361, -32'd915, 32'd7433, -32'd1566},
{-32'd2032, -32'd5230, -32'd8122, -32'd13403},
{32'd5084, 32'd1443, 32'd6582, 32'd5078},
{32'd10798, 32'd8769, 32'd2740, 32'd6209},
{-32'd992, 32'd3480, 32'd11558, 32'd5709},
{32'd3097, -32'd6986, 32'd5460, 32'd6255},
{-32'd6734, 32'd10177, 32'd6490, -32'd13757},
{-32'd4073, -32'd7438, 32'd1738, 32'd3205},
{32'd4075, 32'd12792, 32'd5911, -32'd6953},
{32'd8196, 32'd6512, 32'd510, -32'd2922},
{32'd9615, 32'd8678, -32'd13883, 32'd11492},
{-32'd12779, -32'd15592, 32'd11208, -32'd3876},
{32'd15173, 32'd1005, 32'd16316, 32'd2166},
{-32'd14129, -32'd19218, -32'd73, -32'd4398},
{32'd2059, 32'd3222, 32'd2218, -32'd598},
{-32'd7849, -32'd755, -32'd3629, 32'd2736},
{32'd1404, 32'd262, 32'd15762, 32'd7348},
{-32'd6098, 32'd2441, -32'd3280, -32'd1562},
{32'd2595, -32'd8145, -32'd2191, 32'd6429},
{32'd7551, -32'd12269, 32'd4245, 32'd7585},
{32'd13742, -32'd7550, -32'd9008, 32'd1172},
{-32'd3073, -32'd5698, 32'd759, 32'd4333},
{-32'd5021, -32'd4065, 32'd3175, 32'd5253},
{-32'd10726, -32'd7179, 32'd3280, 32'd6003},
{32'd8993, -32'd9283, 32'd4679, -32'd1323},
{-32'd9082, 32'd7334, 32'd1400, 32'd9851},
{-32'd105, -32'd9823, -32'd14742, 32'd4164},
{32'd10509, 32'd24343, 32'd652, -32'd6936},
{32'd1562, 32'd6767, 32'd5380, 32'd3940},
{-32'd6419, -32'd2478, -32'd1492, 32'd1473},
{-32'd5498, 32'd5610, 32'd11138, 32'd14463},
{-32'd10522, -32'd9863, 32'd5469, -32'd4412},
{32'd886, 32'd19244, -32'd4833, -32'd3051},
{-32'd112, -32'd9789, 32'd11324, 32'd2764},
{32'd15902, 32'd4393, 32'd1218, -32'd4594},
{32'd10342, -32'd14872, 32'd4318, -32'd14865},
{-32'd8323, 32'd7584, -32'd4328, 32'd2867},
{-32'd675, -32'd4520, 32'd3672, -32'd10717},
{32'd733, 32'd14914, 32'd11314, 32'd1696},
{32'd7118, -32'd8125, -32'd2819, -32'd1467},
{32'd1913, -32'd2567, -32'd13942, 32'd1800},
{32'd12349, 32'd1469, 32'd1368, -32'd17848},
{-32'd7206, -32'd3958, -32'd1780, -32'd13769},
{-32'd7878, -32'd9284, 32'd14890, 32'd5519},
{-32'd11847, -32'd12787, -32'd6668, -32'd5894},
{32'd15362, 32'd295, -32'd11318, 32'd4444},
{-32'd1145, -32'd1165, 32'd3881, -32'd11075},
{-32'd6643, -32'd5951, 32'd3158, -32'd2709},
{32'd8758, 32'd4702, 32'd9454, -32'd399},
{-32'd2846, -32'd16580, -32'd447, 32'd4364},
{-32'd5602, -32'd14853, -32'd10734, -32'd9075},
{32'd23944, 32'd6650, 32'd3869, -32'd3962},
{-32'd13749, 32'd2242, 32'd9822, -32'd4237},
{-32'd1803, -32'd8172, 32'd5796, 32'd10705},
{32'd210, 32'd1989, -32'd3818, -32'd2357},
{-32'd5247, -32'd9414, -32'd2041, 32'd1545},
{32'd10224, 32'd11540, 32'd784, 32'd7671},
{-32'd13353, 32'd6345, -32'd13343, 32'd2019},
{-32'd4454, -32'd16696, -32'd10669, 32'd11687},
{32'd8048, -32'd3879, -32'd3122, 32'd1217},
{32'd1990, -32'd6551, 32'd5481, 32'd8081},
{-32'd6467, 32'd1767, 32'd7373, 32'd6316},
{-32'd1912, -32'd5031, 32'd2311, 32'd3913},
{32'd10658, 32'd4998, -32'd5824, 32'd7845},
{-32'd2515, 32'd17450, 32'd3702, 32'd113},
{32'd11554, 32'd6163, -32'd3947, -32'd2482},
{32'd4975, -32'd10969, 32'd2778, 32'd15287},
{-32'd3777, 32'd13168, 32'd12379, 32'd10312},
{32'd2528, 32'd2106, -32'd250, 32'd1251},
{32'd9653, 32'd1164, -32'd9019, -32'd943},
{-32'd5926, 32'd20568, 32'd2521, -32'd280},
{-32'd5807, 32'd11796, -32'd1094, -32'd1356},
{-32'd14404, 32'd9388, -32'd2411, -32'd346},
{-32'd7999, -32'd3374, -32'd2235, 32'd7419},
{32'd9804, 32'd31751, -32'd7768, -32'd6378},
{-32'd2727, -32'd3317, 32'd4743, -32'd9285},
{-32'd1550, 32'd863, 32'd7983, 32'd6587},
{-32'd9589, -32'd3125, 32'd10000, 32'd4993},
{32'd8366, 32'd18414, -32'd3255, 32'd331},
{32'd14118, -32'd2362, -32'd10789, -32'd7927},
{-32'd9227, 32'd9058, -32'd2253, 32'd5624},
{-32'd7156, -32'd8171, 32'd8568, 32'd2756},
{32'd2558, -32'd10103, -32'd5265, 32'd2673},
{-32'd4904, 32'd5811, 32'd3931, -32'd8057},
{-32'd13035, -32'd15345, -32'd1850, -32'd1287},
{-32'd1739, 32'd3521, -32'd6786, 32'd1983},
{-32'd1013, 32'd485, 32'd12104, -32'd6210},
{-32'd10168, -32'd6737, -32'd4594, 32'd11305},
{32'd375, -32'd2357, 32'd4498, 32'd6096},
{-32'd10500, -32'd11173, -32'd5111, -32'd617},
{32'd629, -32'd325, 32'd6710, -32'd2174},
{-32'd7472, -32'd3638, -32'd16966, -32'd8566},
{32'd728, -32'd3823, -32'd9334, -32'd3713},
{-32'd6043, 32'd8576, 32'd9616, 32'd4700},
{-32'd2088, 32'd3631, 32'd3316, -32'd7137},
{-32'd2386, 32'd3080, 32'd9215, -32'd6941},
{32'd720, 32'd8831, 32'd12738, 32'd1885},
{-32'd17393, -32'd8180, 32'd4169, 32'd946},
{32'd2593, 32'd6924, 32'd2473, -32'd5977},
{-32'd2060, 32'd16597, 32'd1867, -32'd4687},
{-32'd12226, 32'd6402, 32'd2452, -32'd3753},
{32'd7427, -32'd3091, -32'd13368, -32'd1935},
{32'd6269, -32'd4237, 32'd13980, 32'd5952},
{32'd3738, 32'd2655, 32'd948, -32'd1690},
{32'd6037, 32'd9102, -32'd3106, 32'd984},
{-32'd9804, 32'd3274, -32'd1947, -32'd960},
{-32'd5491, -32'd9121, 32'd8388, -32'd13416},
{32'd2626, -32'd4948, 32'd7159, 32'd10780},
{-32'd613, 32'd9282, -32'd4112, 32'd3319},
{-32'd4290, -32'd13031, -32'd5211, 32'd3732},
{-32'd10672, 32'd7961, -32'd3415, -32'd4880},
{32'd4056, 32'd4812, -32'd763, 32'd320},
{32'd18615, 32'd10281, 32'd9955, 32'd5257},
{-32'd3842, 32'd10838, 32'd9234, 32'd3825},
{-32'd5385, -32'd15617, -32'd13236, 32'd1923},
{-32'd254, -32'd682, -32'd14890, 32'd4121},
{32'd2298, -32'd2908, 32'd2264, -32'd12500},
{32'd14638, -32'd179, 32'd7229, -32'd6741},
{32'd1221, 32'd1468, 32'd2332, -32'd4890},
{32'd3699, 32'd4990, -32'd3001, -32'd14004},
{32'd229, -32'd4121, 32'd8923, -32'd3578},
{32'd3235, 32'd14177, 32'd7280, -32'd5261},
{32'd4946, -32'd5386, 32'd4428, 32'd1410},
{-32'd12296, -32'd6225, -32'd8799, 32'd1518},
{-32'd1110, 32'd5101, 32'd7631, 32'd3198},
{-32'd4247, 32'd16886, 32'd6197, 32'd2039},
{32'd8430, -32'd17602, -32'd4198, -32'd12883},
{32'd14315, 32'd3753, -32'd2579, -32'd11071},
{-32'd5942, 32'd771, -32'd2671, -32'd8565},
{32'd9662, -32'd178, -32'd396, 32'd4532},
{-32'd4462, -32'd14196, -32'd779, 32'd2659},
{-32'd6894, -32'd2131, 32'd7572, -32'd11748},
{-32'd8324, -32'd11514, -32'd24291, 32'd1390},
{-32'd12177, -32'd6986, -32'd9235, -32'd3137},
{32'd1899, 32'd12006, 32'd1502, -32'd3809},
{-32'd7917, 32'd6171, -32'd4309, 32'd8078},
{32'd12977, -32'd2417, 32'd7095, -32'd13739},
{-32'd1868, -32'd3621, 32'd2696, 32'd2569},
{32'd10050, 32'd2468, -32'd6426, 32'd1890},
{32'd249, 32'd520, -32'd10036, 32'd15409},
{-32'd9949, -32'd9309, 32'd11529, 32'd2805},
{32'd3004, -32'd10475, 32'd1010, 32'd3040},
{32'd10, 32'd1026, 32'd2962, 32'd2360},
{-32'd5945, 32'd152, -32'd8495, -32'd3561},
{32'd112, 32'd5232, 32'd10255, 32'd3294},
{-32'd1249, 32'd8975, 32'd2568, 32'd1820},
{32'd573, -32'd11019, 32'd4659, 32'd7881},
{32'd5883, -32'd9780, 32'd2031, 32'd8367},
{32'd17967, 32'd80, 32'd7142, 32'd3139},
{-32'd2875, -32'd19918, -32'd2636, 32'd10278},
{-32'd9204, 32'd8734, 32'd13284, 32'd5882},
{32'd4989, 32'd2358, 32'd10077, -32'd3376},
{-32'd8867, 32'd1930, -32'd10159, 32'd11389},
{32'd8638, -32'd1428, 32'd118, -32'd4312},
{-32'd602, 32'd5430, -32'd3675, -32'd5770},
{32'd1629, 32'd19586, -32'd6474, 32'd7103},
{32'd10762, -32'd9573, -32'd3614, -32'd12056},
{32'd14728, 32'd1859, -32'd1, -32'd6710},
{32'd2305, -32'd4927, 32'd12646, -32'd2607},
{32'd9916, -32'd11686, 32'd6987, -32'd8166},
{32'd3297, -32'd13042, 32'd1071, -32'd7990},
{-32'd1028, 32'd3467, 32'd8751, 32'd6622},
{-32'd1691, -32'd2604, 32'd10257, -32'd4645},
{-32'd7517, 32'd7263, 32'd15627, -32'd6142},
{32'd9590, -32'd9805, -32'd8061, -32'd8445},
{32'd528, -32'd10800, 32'd6765, 32'd7218},
{32'd2805, 32'd16173, 32'd9434, -32'd8251},
{32'd7496, -32'd5778, -32'd952, 32'd6431},
{-32'd11678, 32'd2093, -32'd8796, -32'd49},
{-32'd11901, 32'd982, 32'd7991, -32'd5872},
{-32'd12275, -32'd7833, -32'd6457, -32'd5331},
{32'd1782, -32'd5403, -32'd3102, -32'd8876},
{32'd7333, 32'd3759, -32'd3978, -32'd2268},
{32'd1682, 32'd1014, 32'd1892, -32'd1437},
{32'd12663, -32'd14692, -32'd1997, 32'd6381},
{-32'd428, -32'd6545, 32'd1441, 32'd6590},
{32'd4660, 32'd2826, -32'd2439, 32'd4996},
{32'd12176, -32'd9461, -32'd177, 32'd3000},
{-32'd2338, -32'd18574, 32'd336, 32'd4004},
{-32'd13532, 32'd9422, 32'd4313, 32'd5132},
{-32'd8488, -32'd9713, -32'd8193, -32'd13999},
{32'd6488, -32'd2912, 32'd8501, 32'd3951},
{32'd7777, -32'd10007, 32'd2264, -32'd16},
{-32'd2158, 32'd1252, 32'd5553, 32'd2285},
{-32'd1726, -32'd4732, -32'd669, 32'd10057},
{-32'd2690, 32'd6461, 32'd6438, -32'd1008},
{32'd15474, -32'd8011, -32'd6149, -32'd8677},
{32'd7470, 32'd1299, -32'd2392, -32'd1832},
{32'd3287, -32'd2788, 32'd4009, 32'd1524},
{-32'd6768, -32'd2088, -32'd5682, -32'd6340},
{32'd8607, -32'd11020, -32'd3002, -32'd12223},
{-32'd7382, -32'd5808, -32'd7695, 32'd812},
{-32'd5283, -32'd3751, -32'd705, -32'd80},
{32'd16712, -32'd4789, -32'd9438, 32'd1965},
{-32'd5382, 32'd12762, -32'd882, -32'd1161},
{32'd7204, -32'd2750, 32'd8621, 32'd10628},
{-32'd16035, -32'd1217, -32'd2305, 32'd191},
{32'd12976, -32'd2857, -32'd9545, 32'd2063},
{32'd6854, 32'd13711, -32'd13842, -32'd2242},
{-32'd697, 32'd10373, 32'd4890, 32'd1392},
{-32'd11354, -32'd5111, -32'd3914, 32'd7285},
{-32'd3025, 32'd16076, -32'd7378, -32'd1030},
{-32'd1747, 32'd8076, -32'd14382, -32'd6834},
{32'd6620, 32'd2983, -32'd4233, -32'd531},
{-32'd8112, -32'd9738, 32'd12746, 32'd8189},
{-32'd1667, -32'd2821, -32'd15479, -32'd9439},
{32'd12580, -32'd14893, -32'd5943, -32'd3854},
{-32'd9795, -32'd10935, 32'd5806, 32'd12570},
{32'd2159, 32'd13454, 32'd2940, -32'd333},
{32'd2088, 32'd10216, -32'd5221, -32'd9793},
{32'd5893, 32'd11635, -32'd3490, -32'd6058},
{32'd5062, -32'd9589, 32'd7687, -32'd6112},
{-32'd922, -32'd8000, -32'd7083, 32'd787},
{32'd6498, 32'd1341, 32'd309, -32'd2333},
{-32'd11352, -32'd4827, -32'd6289, 32'd8140},
{-32'd13366, -32'd7374, -32'd2091, -32'd1347},
{32'd1590, -32'd4828, -32'd5357, 32'd7107},
{-32'd2161, 32'd11491, -32'd7172, -32'd35},
{32'd6200, 32'd2964, 32'd6051, 32'd4577},
{32'd7579, 32'd15795, 32'd5025, -32'd5328},
{-32'd6468, 32'd2994, 32'd10699, -32'd7188},
{32'd6004, -32'd2379, -32'd4539, -32'd488},
{32'd5309, 32'd11792, 32'd12288, 32'd2209},
{-32'd9195, -32'd7049, -32'd12857, -32'd8289},
{32'd1785, -32'd7245, -32'd6465, 32'd8188},
{32'd3828, -32'd7888, -32'd2515, 32'd5309},
{32'd11224, -32'd1068, 32'd10256, 32'd8004},
{-32'd19088, -32'd4074, -32'd656, -32'd6946},
{32'd5916, -32'd10849, 32'd3171, 32'd2304},
{32'd16357, 32'd12692, 32'd497, -32'd6441},
{32'd3293, -32'd11561, -32'd16127, -32'd9011},
{-32'd7491, -32'd366, -32'd2894, -32'd2996},
{32'd4420, 32'd8234, -32'd7341, -32'd3720},
{-32'd10574, 32'd6170, -32'd271, -32'd9648},
{32'd4265, -32'd13650, -32'd954, -32'd6268},
{-32'd4556, 32'd4307, -32'd3263, -32'd2697},
{-32'd3470, -32'd631, 32'd6476, -32'd2270},
{-32'd4507, 32'd5138, -32'd8655, -32'd4335},
{-32'd12254, 32'd389, -32'd2918, -32'd1255},
{-32'd15332, -32'd10474, -32'd5180, -32'd2811},
{32'd3460, 32'd4795, 32'd2320, -32'd8329},
{-32'd1704, 32'd439, -32'd4182, 32'd1184},
{-32'd14132, -32'd6721, 32'd288, 32'd6016},
{-32'd9957, -32'd16270, -32'd9258, 32'd2697},
{32'd17169, 32'd8007, -32'd1630, -32'd1773},
{32'd790, -32'd813, 32'd3773, 32'd4865},
{-32'd9910, 32'd17171, -32'd8010, -32'd17022},
{32'd3635, -32'd8135, -32'd3518, -32'd10140},
{-32'd5435, 32'd1444, -32'd3185, -32'd220},
{32'd3639, 32'd16302, 32'd11259, 32'd8974},
{-32'd2349, -32'd11890, -32'd5373, 32'd8010},
{-32'd1575, -32'd2642, 32'd7923, -32'd15454},
{-32'd5375, 32'd7843, -32'd4234, -32'd3205},
{32'd7203, 32'd2785, 32'd9027, 32'd17424},
{-32'd7122, -32'd5212, 32'd3632, 32'd4982},
{32'd5907, -32'd12749, -32'd6949, -32'd18589},
{32'd2998, 32'd2759, 32'd13237, 32'd14253},
{-32'd3126, -32'd12176, -32'd6107, -32'd4065},
{-32'd3331, -32'd12301, 32'd1594, 32'd1188},
{-32'd4077, 32'd14848, 32'd1844, -32'd16277},
{-32'd534, -32'd228, 32'd1095, 32'd815},
{-32'd3813, 32'd1358, 32'd9176, -32'd1051},
{-32'd12670, 32'd2556, -32'd882, -32'd9951},
{-32'd3520, 32'd10210, -32'd51, 32'd791},
{-32'd3953, -32'd969, 32'd65, -32'd7852},
{-32'd14024, -32'd1243, 32'd5375, -32'd2507},
{-32'd6284, 32'd10017, 32'd2360, -32'd3985},
{32'd14225, -32'd3746, -32'd1586, -32'd4461},
{-32'd6458, -32'd7752, -32'd3193, -32'd9032},
{-32'd9487, -32'd4808, -32'd1346, 32'd13688},
{32'd5313, 32'd9528, 32'd145, 32'd8766},
{32'd6937, 32'd2030, -32'd832, -32'd12467},
{-32'd6964, 32'd11382, 32'd8912, 32'd4266},
{-32'd7199, -32'd410, -32'd10028, -32'd2391},
{-32'd4489, 32'd12747, 32'd19339, 32'd7914},
{-32'd2162, -32'd8546, -32'd4094, -32'd4840},
{32'd11006, 32'd6267, 32'd306, -32'd2098},
{-32'd2882, -32'd6025, -32'd4439, -32'd11631},
{-32'd11230, -32'd1946, -32'd135, 32'd3496},
{32'd7090, -32'd1789, 32'd4002, 32'd9258},
{32'd5242, 32'd3499, 32'd10459, -32'd4642},
{32'd7241, 32'd13629, 32'd589, -32'd2064},
{-32'd6316, 32'd17544, -32'd2566, -32'd5257},
{32'd2995, 32'd11892, -32'd7249, -32'd17013},
{32'd12356, -32'd2208, -32'd4153, 32'd7677},
{-32'd13440, -32'd9501, -32'd1329, 32'd11477},
{32'd1629, 32'd10619, -32'd2468, 32'd6270},
{-32'd8194, 32'd8549, -32'd3332, -32'd9795},
{-32'd1556, 32'd2048, 32'd9473, -32'd15912},
{32'd2362, -32'd8860, -32'd4189, -32'd3124},
{-32'd2357, -32'd24991, -32'd3348, 32'd10884},
{32'd9282, 32'd7911, -32'd9511, 32'd779},
{-32'd1198, -32'd19620, -32'd7285, -32'd3836},
{32'd5770, -32'd1893, -32'd926, -32'd5623},
{-32'd14791, 32'd2749, -32'd21732, -32'd7329},
{-32'd1260, 32'd7906, 32'd4064, -32'd2537},
{-32'd6085, -32'd3937, -32'd3957, -32'd10227},
{32'd11250, 32'd6932, 32'd2955, 32'd6453},
{32'd11321, -32'd6331, 32'd9321, 32'd1204},
{-32'd8185, -32'd7073, 32'd1117, 32'd282}
},
{{-32'd11297, 32'd8754, -32'd1884, -32'd8032},
{-32'd1480, -32'd6348, -32'd4903, -32'd919},
{32'd1845, -32'd2091, -32'd788, 32'd7725},
{-32'd1860, 32'd6097, -32'd700, -32'd921},
{-32'd4063, 32'd10079, 32'd580, -32'd1440},
{-32'd6127, 32'd3598, 32'd7602, 32'd5570},
{-32'd1847, 32'd8441, 32'd6578, -32'd12691},
{-32'd8622, -32'd8581, -32'd2292, -32'd9405},
{-32'd14347, -32'd811, 32'd9189, 32'd5761},
{32'd5497, 32'd22430, 32'd5437, 32'd2273},
{-32'd1839, -32'd508, 32'd4066, 32'd3349},
{32'd8173, -32'd2314, -32'd1354, -32'd974},
{-32'd5976, 32'd3596, 32'd7792, 32'd1335},
{32'd13, -32'd2127, -32'd9850, 32'd12878},
{-32'd6505, -32'd7109, 32'd2689, -32'd14978},
{-32'd17964, -32'd5699, -32'd6376, -32'd7607},
{-32'd924, -32'd6572, 32'd4744, 32'd2760},
{-32'd8110, 32'd1180, -32'd6660, 32'd20151},
{32'd1749, 32'd6160, 32'd2483, 32'd5537},
{32'd5991, 32'd1723, -32'd6801, -32'd4628},
{32'd2885, -32'd9739, 32'd3733, -32'd1396},
{-32'd5386, -32'd2060, -32'd10566, -32'd3122},
{-32'd3414, -32'd1998, 32'd9916, -32'd3101},
{32'd3059, -32'd11561, -32'd486, 32'd2007},
{32'd10508, -32'd1009, 32'd806, 32'd8969},
{-32'd10671, 32'd3481, -32'd9314, -32'd826},
{32'd3989, -32'd7625, 32'd2116, -32'd6299},
{32'd11974, 32'd7988, 32'd15061, 32'd5033},
{32'd3397, 32'd9239, 32'd2228, 32'd5499},
{-32'd599, -32'd4079, 32'd4814, 32'd12638},
{32'd3242, -32'd1006, 32'd2655, 32'd4554},
{-32'd3554, 32'd53, -32'd4885, -32'd4673},
{32'd1995, 32'd11078, 32'd7427, 32'd908},
{32'd2475, 32'd3007, -32'd9160, 32'd4589},
{32'd702, 32'd10249, 32'd8185, -32'd662},
{-32'd4170, -32'd6246, -32'd5542, -32'd6504},
{32'd927, 32'd14300, 32'd2213, -32'd3638},
{-32'd13006, -32'd8146, -32'd5775, 32'd1257},
{32'd2866, -32'd5459, 32'd825, -32'd73},
{32'd4354, 32'd429, -32'd1635, -32'd4787},
{-32'd4925, -32'd5940, -32'd2401, -32'd5135},
{32'd4652, 32'd6171, -32'd7227, 32'd2890},
{32'd10907, -32'd4714, -32'd2569, 32'd5928},
{-32'd2095, 32'd9690, -32'd5799, -32'd1625},
{-32'd5349, -32'd5684, 32'd2662, -32'd5111},
{32'd9522, 32'd9937, -32'd10376, 32'd9055},
{-32'd3939, 32'd240, 32'd1869, -32'd7566},
{32'd163, -32'd4581, -32'd6219, 32'd4507},
{-32'd783, -32'd2876, 32'd13183, 32'd376},
{-32'd3541, 32'd147, 32'd4622, -32'd4751},
{-32'd819, -32'd1528, -32'd3948, 32'd1436},
{32'd5798, -32'd10085, -32'd7747, -32'd7431},
{32'd5101, -32'd5691, 32'd3434, -32'd8349},
{-32'd1839, -32'd5249, 32'd1433, -32'd1559},
{-32'd7788, 32'd9154, 32'd11080, 32'd7355},
{-32'd1096, 32'd3178, -32'd11849, 32'd3708},
{-32'd3180, -32'd1187, -32'd1679, 32'd7970},
{-32'd2546, 32'd188, -32'd1583, -32'd8527},
{32'd536, -32'd9288, -32'd4720, 32'd5499},
{32'd1713, -32'd5321, 32'd2163, 32'd4872},
{32'd3278, -32'd3805, -32'd7467, -32'd10376},
{-32'd4489, -32'd2822, -32'd10651, 32'd8011},
{-32'd411, -32'd16112, -32'd5374, -32'd1454},
{-32'd3811, 32'd257, -32'd961, -32'd7088},
{32'd825, 32'd5912, -32'd3450, -32'd7528},
{32'd4411, 32'd10710, 32'd4793, 32'd1322},
{32'd5731, -32'd7268, 32'd7473, -32'd3243},
{-32'd2353, -32'd5923, 32'd2182, -32'd2559},
{32'd523, -32'd666, -32'd3935, 32'd8043},
{32'd3602, -32'd4016, 32'd1321, -32'd7846},
{-32'd5573, 32'd3835, -32'd1326, -32'd3405},
{32'd234, -32'd7681, -32'd1598, 32'd2501},
{-32'd9958, 32'd1268, 32'd5944, 32'd792},
{-32'd5653, -32'd1480, -32'd3081, 32'd3780},
{32'd1636, 32'd506, -32'd2047, 32'd2894},
{32'd2479, -32'd7592, -32'd9112, -32'd3169},
{-32'd1178, -32'd3553, -32'd8205, 32'd9301},
{32'd4831, -32'd4714, -32'd2596, 32'd11890},
{32'd8565, 32'd2037, 32'd3767, -32'd972},
{-32'd3560, -32'd4066, -32'd10648, -32'd1491},
{-32'd552, 32'd9135, 32'd6965, -32'd14607},
{32'd7099, 32'd7297, 32'd1691, -32'd1731},
{-32'd4734, 32'd948, -32'd170, -32'd3239},
{-32'd3088, -32'd3912, 32'd150, 32'd1829},
{-32'd4104, 32'd4411, -32'd7846, 32'd5047},
{32'd8116, 32'd5603, 32'd2294, 32'd4070},
{32'd1992, 32'd8638, -32'd3797, -32'd3910},
{-32'd9075, -32'd21875, -32'd5184, -32'd7439},
{32'd5346, 32'd4957, -32'd6812, 32'd6330},
{32'd5575, -32'd14175, -32'd7806, -32'd5675},
{-32'd1494, 32'd13116, 32'd4784, 32'd2812},
{32'd1309, -32'd2587, 32'd1598, -32'd2660},
{-32'd1160, 32'd10476, 32'd4307, 32'd3632},
{32'd3598, 32'd453, -32'd1776, 32'd4263},
{-32'd2011, 32'd534, -32'd2501, 32'd6695},
{-32'd1450, -32'd113, -32'd3795, -32'd8291},
{32'd4000, 32'd13791, 32'd6138, -32'd2023},
{-32'd9429, -32'd930, 32'd8079, 32'd1238},
{32'd3417, -32'd5775, -32'd3506, -32'd11772},
{32'd581, 32'd9549, -32'd2257, -32'd3450},
{32'd4546, -32'd7922, -32'd4402, 32'd1415},
{-32'd662, -32'd2686, -32'd433, 32'd1333},
{32'd3963, 32'd8960, 32'd7768, 32'd2568},
{32'd3400, 32'd2398, 32'd4512, -32'd11953},
{32'd8773, -32'd10313, 32'd10694, -32'd2503},
{-32'd8306, -32'd26, 32'd437, -32'd9916},
{-32'd8441, -32'd2433, 32'd3283, 32'd4006},
{-32'd7568, -32'd5028, -32'd932, 32'd2749},
{32'd5931, 32'd18212, 32'd10691, 32'd1167},
{-32'd1479, -32'd8136, 32'd2651, -32'd10203},
{32'd3709, -32'd3103, -32'd6285, -32'd6015},
{32'd2983, -32'd689, -32'd4147, -32'd2386},
{32'd3183, 32'd19003, 32'd9701, -32'd1825},
{32'd5429, 32'd10120, -32'd6076, -32'd251},
{-32'd11258, 32'd2863, -32'd5751, -32'd7190},
{32'd5818, -32'd9473, 32'd4443, -32'd1367},
{32'd1299, -32'd301, 32'd2696, 32'd835},
{32'd3347, 32'd419, 32'd3900, 32'd3875},
{-32'd5907, -32'd7338, 32'd1121, -32'd10921},
{32'd8856, 32'd9951, 32'd6584, -32'd3130},
{32'd1883, 32'd1909, -32'd3025, 32'd877},
{32'd13300, -32'd8120, 32'd3121, 32'd7094},
{32'd2788, -32'd7079, -32'd4746, -32'd3920},
{32'd1761, -32'd5025, 32'd3742, -32'd530},
{32'd241, 32'd8441, 32'd2120, -32'd2655},
{-32'd3354, 32'd5651, 32'd7053, 32'd8009},
{-32'd982, -32'd9486, -32'd1672, 32'd2038},
{32'd9705, -32'd15235, -32'd6483, -32'd5188},
{-32'd6499, 32'd704, -32'd2726, -32'd6300},
{32'd1586, -32'd1029, 32'd5026, 32'd1654},
{-32'd1779, 32'd2717, -32'd92, -32'd4667},
{-32'd6907, -32'd6332, 32'd572, -32'd721},
{32'd1779, -32'd1577, 32'd5182, 32'd766},
{32'd3058, 32'd3579, -32'd4046, -32'd5413},
{-32'd264, -32'd9293, 32'd1380, 32'd2585},
{32'd4639, 32'd2002, -32'd3523, 32'd1397},
{-32'd1025, 32'd3338, 32'd1060, 32'd8312},
{32'd1093, -32'd2097, -32'd2183, -32'd10193},
{32'd5111, -32'd11014, 32'd10928, 32'd2590},
{32'd1944, -32'd14779, -32'd3369, 32'd1002},
{-32'd518, 32'd2274, 32'd9398, 32'd626},
{-32'd2278, -32'd4611, -32'd2143, -32'd7533},
{-32'd5535, -32'd6653, 32'd2703, -32'd3028},
{-32'd14400, 32'd4860, 32'd2841, -32'd10455},
{32'd12347, 32'd12059, -32'd4028, 32'd5210},
{-32'd648, 32'd610, -32'd2219, -32'd8170},
{32'd3040, -32'd4865, 32'd6890, 32'd12554},
{-32'd8142, -32'd560, -32'd5192, -32'd2755},
{32'd4170, -32'd13481, -32'd3843, -32'd12410},
{-32'd2014, 32'd2011, -32'd206, -32'd2487},
{32'd4991, -32'd5872, 32'd2899, 32'd673},
{32'd4513, 32'd2341, 32'd13839, -32'd4577},
{-32'd4994, -32'd955, 32'd4239, -32'd2550},
{32'd4763, -32'd2048, -32'd12796, 32'd1593},
{32'd192, -32'd7339, 32'd6026, -32'd1670},
{-32'd4062, 32'd8296, 32'd4189, -32'd6571},
{32'd2053, -32'd5689, 32'd1797, 32'd806},
{-32'd4045, -32'd3787, 32'd2465, 32'd14138},
{32'd6772, -32'd2211, -32'd344, -32'd7922},
{-32'd6499, -32'd1276, -32'd1364, 32'd4464},
{-32'd11398, 32'd3527, -32'd5862, 32'd4515},
{32'd6505, 32'd4485, 32'd2162, 32'd848},
{32'd4845, -32'd12083, 32'd4320, -32'd4444},
{32'd1178, 32'd36, 32'd10562, -32'd3431},
{32'd1463, -32'd4915, 32'd6020, 32'd3300},
{32'd7338, -32'd663, -32'd1155, 32'd603},
{-32'd6629, 32'd6229, -32'd2903, 32'd1155},
{32'd2627, -32'd15948, -32'd7063, -32'd1184},
{-32'd2704, 32'd807, -32'd6868, 32'd6440},
{-32'd4550, -32'd12877, -32'd3694, 32'd6533},
{32'd341, 32'd1544, -32'd5789, 32'd4794},
{-32'd2020, 32'd5294, -32'd763, -32'd3793},
{32'd2059, 32'd9259, 32'd6989, 32'd224},
{-32'd3196, 32'd4957, -32'd13027, 32'd537},
{32'd11861, -32'd5924, 32'd5730, -32'd6266},
{32'd6680, 32'd10719, 32'd825, 32'd11717},
{-32'd661, 32'd3296, 32'd12398, 32'd3963},
{-32'd2919, -32'd4603, 32'd4536, -32'd529},
{-32'd13168, 32'd9656, 32'd7066, -32'd10455},
{-32'd2522, -32'd7279, -32'd970, -32'd7432},
{-32'd5285, 32'd538, -32'd4089, -32'd4616},
{-32'd6693, -32'd1337, 32'd4628, -32'd8560},
{-32'd5902, -32'd8820, -32'd1385, -32'd7123},
{-32'd8090, 32'd9592, -32'd5821, -32'd10559},
{32'd1223, 32'd14691, 32'd10922, 32'd7404},
{-32'd2128, -32'd4223, 32'd7345, -32'd519},
{32'd1698, 32'd5004, 32'd5739, -32'd7255},
{-32'd8554, -32'd1541, 32'd1955, -32'd10036},
{-32'd7042, 32'd1000, -32'd5452, -32'd1454},
{32'd7057, 32'd5773, -32'd9205, -32'd3715},
{-32'd8717, -32'd3252, 32'd2484, -32'd6204},
{32'd4156, -32'd8998, -32'd5820, 32'd129},
{-32'd2831, -32'd7110, 32'd928, 32'd1357},
{32'd3313, -32'd2230, -32'd272, -32'd1593},
{-32'd6484, -32'd6760, 32'd3779, -32'd6939},
{-32'd3354, 32'd5738, 32'd12795, -32'd436},
{-32'd9429, -32'd10899, 32'd5888, -32'd12333},
{32'd8431, -32'd3161, -32'd2480, 32'd7598},
{-32'd5103, -32'd2454, -32'd145, -32'd6854},
{-32'd3640, -32'd670, 32'd7136, 32'd101},
{-32'd3903, -32'd8456, -32'd3165, -32'd1191},
{-32'd4158, 32'd3395, 32'd11051, -32'd5896},
{32'd2822, -32'd834, -32'd947, -32'd23051},
{32'd4996, 32'd7379, 32'd4374, -32'd6681},
{32'd1765, -32'd7080, -32'd13224, 32'd3440},
{32'd12692, -32'd5788, 32'd3512, -32'd4743},
{-32'd9200, -32'd3507, 32'd3441, -32'd5412},
{32'd5975, 32'd10155, 32'd5101, -32'd9396},
{-32'd8424, 32'd2480, 32'd646, -32'd7230},
{32'd4147, -32'd4995, -32'd6093, 32'd5274},
{-32'd1449, -32'd2008, -32'd5930, -32'd5662},
{32'd4259, 32'd2772, -32'd8422, -32'd948},
{-32'd498, -32'd10511, -32'd4509, -32'd2790},
{-32'd5813, -32'd125, -32'd290, -32'd5413},
{-32'd195, 32'd3181, 32'd5686, 32'd3767},
{-32'd1481, -32'd817, 32'd7003, -32'd4058},
{-32'd10899, 32'd164, -32'd5705, -32'd1317},
{-32'd6627, -32'd6478, 32'd10941, -32'd4440},
{32'd8105, 32'd613, -32'd875, 32'd8477},
{-32'd2768, -32'd14080, -32'd347, -32'd1485},
{-32'd178, -32'd727, -32'd7624, -32'd3586},
{-32'd1342, 32'd717, 32'd7226, -32'd2197},
{-32'd1495, 32'd9651, 32'd11880, -32'd8591},
{32'd3930, -32'd566, 32'd5763, 32'd7719},
{-32'd4939, 32'd4980, -32'd2032, -32'd1359},
{-32'd3080, 32'd5309, -32'd6566, -32'd6310},
{-32'd713, -32'd9239, -32'd3987, -32'd1589},
{32'd4466, -32'd9637, 32'd877, 32'd1080},
{-32'd1347, -32'd4635, 32'd2733, -32'd2266},
{-32'd12, -32'd11456, -32'd11683, -32'd4080},
{-32'd5761, -32'd3713, 32'd8261, 32'd4070},
{32'd3468, 32'd6821, -32'd3480, 32'd8849},
{-32'd7203, -32'd5920, -32'd4268, -32'd2698},
{-32'd4061, 32'd6685, 32'd7697, -32'd33},
{-32'd1552, 32'd3136, -32'd15894, 32'd4455},
{-32'd1791, -32'd2726, -32'd8492, 32'd2624},
{32'd2338, 32'd10656, 32'd4710, -32'd1711},
{-32'd1352, 32'd8207, 32'd4249, 32'd3086},
{32'd2399, 32'd579, 32'd6087, 32'd2486},
{32'd2373, -32'd5756, -32'd3122, 32'd3423},
{-32'd1528, -32'd7911, -32'd3228, 32'd3403},
{32'd2300, -32'd6452, -32'd3974, 32'd1536},
{-32'd7342, -32'd12358, 32'd481, -32'd1546},
{32'd259, 32'd9540, -32'd17171, -32'd5371},
{32'd1041, 32'd18913, 32'd6878, 32'd1799},
{32'd7363, -32'd1963, 32'd8559, 32'd372},
{-32'd7883, -32'd7099, 32'd719, -32'd12474},
{32'd3002, -32'd6304, 32'd1733, 32'd12429},
{-32'd7773, -32'd4653, -32'd4014, -32'd495},
{-32'd4873, -32'd3519, -32'd10290, 32'd488},
{-32'd6707, 32'd2346, 32'd981, 32'd8638},
{32'd2613, 32'd5154, 32'd5932, 32'd8202},
{32'd1683, 32'd5168, -32'd6549, 32'd1320},
{-32'd13522, 32'd6603, -32'd2418, -32'd2262},
{-32'd9855, -32'd10626, 32'd5713, -32'd6598},
{-32'd576, 32'd397, -32'd7696, -32'd3556},
{-32'd1125, 32'd5024, 32'd5531, 32'd2644},
{32'd4884, 32'd6763, 32'd1184, -32'd9448},
{-32'd10203, 32'd4530, -32'd1482, -32'd3851},
{-32'd926, 32'd136, -32'd15107, 32'd10049},
{-32'd11488, 32'd7223, 32'd7592, 32'd3893},
{32'd6315, -32'd150, -32'd11664, 32'd4964},
{32'd2980, 32'd345, -32'd13692, -32'd409},
{32'd3391, -32'd3361, -32'd6449, -32'd7645},
{32'd1375, 32'd11535, 32'd9290, -32'd4993},
{-32'd3642, -32'd6218, -32'd8234, -32'd5304},
{32'd4545, 32'd9198, 32'd5581, 32'd2684},
{-32'd4176, -32'd10628, 32'd239, 32'd4140},
{-32'd1528, -32'd3323, 32'd1445, 32'd4676},
{32'd3875, -32'd4577, -32'd6290, -32'd4619},
{-32'd468, -32'd2273, 32'd7057, 32'd6361},
{-32'd3590, 32'd1261, 32'd4348, -32'd5794},
{32'd1967, -32'd10273, -32'd2409, -32'd7343},
{-32'd5426, -32'd8217, 32'd4843, 32'd5310},
{-32'd12400, -32'd7894, -32'd15574, 32'd6874},
{32'd5186, -32'd4398, 32'd510, -32'd248},
{32'd5217, 32'd17604, 32'd3770, 32'd2050},
{32'd4251, -32'd2400, 32'd4065, 32'd1543},
{-32'd3485, -32'd17691, -32'd4365, -32'd947},
{32'd1512, -32'd2615, -32'd2526, -32'd4471},
{-32'd1604, 32'd1517, 32'd1252, 32'd816},
{-32'd2802, 32'd713, 32'd1903, -32'd9600},
{-32'd5872, -32'd2218, -32'd3803, 32'd8869},
{32'd7435, -32'd5920, -32'd7645, -32'd3479},
{32'd1865, -32'd5918, 32'd510, 32'd6443},
{-32'd647, -32'd9083, -32'd4302, -32'd8170},
{32'd5172, 32'd5923, 32'd9450, 32'd538},
{32'd8259, -32'd10172, 32'd4225, -32'd6465},
{32'd1819, 32'd5317, -32'd6482, -32'd4388},
{32'd2943, 32'd14, -32'd11187, 32'd2841},
{32'd1767, -32'd1788, 32'd5550, -32'd6431},
{32'd5077, 32'd9361, 32'd1599, 32'd7819},
{-32'd5958, -32'd11161, 32'd3010, -32'd11348},
{32'd515, -32'd314, 32'd2244, 32'd3959},
{32'd3278, -32'd12658, -32'd5983, -32'd4864},
{-32'd3721, -32'd11144, -32'd2661, -32'd349},
{-32'd612, 32'd992, 32'd2785, 32'd4300},
{32'd1407, -32'd1358, 32'd354, -32'd145},
{-32'd2103, 32'd2650, 32'd1053, 32'd3807},
{-32'd8530, 32'd6641, -32'd9360, -32'd11735}
},
{{32'd8171, 32'd7429, 32'd3460, -32'd5668},
{32'd1373, 32'd905, -32'd2834, -32'd3270},
{-32'd3129, 32'd8544, 32'd5284, 32'd1391},
{-32'd2381, -32'd3057, -32'd3065, -32'd1411},
{-32'd1346, 32'd621, 32'd1586, 32'd2040},
{-32'd5432, -32'd4789, -32'd9394, -32'd1238},
{32'd2611, 32'd5740, 32'd5536, 32'd740},
{-32'd8425, -32'd8672, 32'd187, -32'd2966},
{32'd7007, -32'd7802, -32'd9564, 32'd1778},
{32'd15818, 32'd7469, 32'd6569, 32'd8751},
{32'd5042, 32'd5949, -32'd2489, 32'd3395},
{32'd9711, -32'd1358, -32'd3820, 32'd304},
{-32'd1039, 32'd6392, 32'd1967, -32'd1773},
{32'd3760, -32'd3701, 32'd4479, -32'd5174},
{-32'd3672, -32'd3604, -32'd7585, -32'd337},
{32'd1419, 32'd35, -32'd2030, -32'd1164},
{32'd5344, 32'd10910, -32'd104, 32'd2110},
{-32'd2849, 32'd6444, 32'd10915, 32'd2490},
{32'd7328, -32'd4356, 32'd99, 32'd6432},
{-32'd5152, 32'd2009, 32'd815, -32'd1104},
{32'd398, 32'd2532, 32'd4160, -32'd1669},
{-32'd10836, -32'd8635, 32'd1716, -32'd2205},
{-32'd6991, -32'd737, -32'd2876, 32'd2395},
{-32'd11429, -32'd4737, -32'd1686, -32'd5255},
{32'd2135, 32'd14880, 32'd3973, 32'd5360},
{32'd2924, 32'd6038, 32'd8568, -32'd396},
{-32'd4019, 32'd3447, -32'd1335, -32'd2064},
{32'd303, 32'd4702, -32'd1129, 32'd1781},
{-32'd1405, 32'd121, 32'd8475, 32'd3251},
{32'd1181, -32'd7216, -32'd1547, 32'd4093},
{-32'd1614, 32'd8665, -32'd1569, -32'd3477},
{-32'd3695, -32'd6597, -32'd602, -32'd6002},
{32'd12272, 32'd1387, -32'd98, 32'd2865},
{-32'd9526, 32'd3257, 32'd2363, -32'd5010},
{32'd6789, 32'd5358, 32'd6248, 32'd3333},
{-32'd7853, 32'd4337, 32'd3079, -32'd1214},
{-32'd2187, -32'd7438, 32'd285, -32'd6376},
{32'd3917, -32'd646, -32'd3738, -32'd405},
{-32'd5170, 32'd2519, -32'd608, 32'd226},
{-32'd10969, 32'd8677, 32'd3500, -32'd3170},
{-32'd3673, 32'd906, 32'd4891, 32'd1210},
{-32'd689, -32'd1800, 32'd4728, -32'd969},
{-32'd118, 32'd6703, 32'd3637, -32'd5743},
{-32'd793, 32'd2295, -32'd186, -32'd4406},
{-32'd1521, -32'd2168, -32'd999, 32'd3300},
{32'd534, -32'd942, -32'd11111, -32'd3050},
{-32'd7766, -32'd599, 32'd1971, 32'd6103},
{-32'd4783, -32'd297, -32'd4213, 32'd2865},
{32'd2963, 32'd5334, -32'd1312, 32'd1364},
{-32'd1383, 32'd1668, -32'd3408, -32'd4051},
{32'd1825, -32'd3166, 32'd709, -32'd5806},
{32'd5487, -32'd13171, 32'd1457, -32'd5046},
{32'd926, -32'd113, -32'd4485, 32'd3696},
{-32'd6304, 32'd7034, 32'd5350, -32'd3821},
{32'd4505, 32'd10077, 32'd2380, 32'd4386},
{32'd4815, 32'd6001, -32'd5408, -32'd5902},
{32'd1257, -32'd4105, 32'd2106, 32'd5308},
{32'd404, -32'd4691, -32'd870, -32'd3891},
{-32'd4503, -32'd3826, -32'd2063, -32'd2885},
{-32'd5630, 32'd5262, -32'd4567, -32'd798},
{-32'd7959, -32'd3286, 32'd624, -32'd2150},
{-32'd1240, 32'd2235, -32'd233, -32'd5683},
{-32'd676, -32'd504, 32'd474, -32'd4445},
{-32'd467, 32'd6892, -32'd1533, 32'd364},
{32'd2054, 32'd3700, -32'd1847, 32'd1870},
{32'd4382, -32'd3562, 32'd4277, 32'd1199},
{-32'd3056, -32'd2062, -32'd569, -32'd1214},
{-32'd4371, 32'd1583, 32'd714, -32'd4175},
{32'd3624, -32'd661, -32'd1931, -32'd1268},
{-32'd1835, -32'd5032, 32'd3738, -32'd2224},
{32'd187, -32'd6430, -32'd2169, 32'd1151},
{32'd1665, -32'd1058, 32'd3994, 32'd1137},
{32'd450, 32'd4480, 32'd2398, -32'd5617},
{32'd45, -32'd4368, -32'd3272, 32'd3383},
{-32'd1170, -32'd312, 32'd755, 32'd6891},
{-32'd6714, 32'd1647, 32'd6796, -32'd5515},
{32'd1828, -32'd3320, -32'd1032, -32'd1381},
{32'd4392, -32'd3015, 32'd2464, 32'd3234},
{32'd3707, -32'd5263, 32'd6992, 32'd238},
{-32'd2706, -32'd2542, 32'd2277, -32'd2554},
{32'd2874, -32'd1907, 32'd785, 32'd5262},
{32'd1631, 32'd6249, 32'd4508, 32'd2099},
{-32'd2861, 32'd1625, 32'd3153, 32'd3523},
{32'd3199, 32'd947, -32'd445, -32'd5299},
{32'd2443, -32'd3283, 32'd4459, -32'd3929},
{32'd1560, 32'd6468, -32'd6688, -32'd2144},
{32'd2728, -32'd3606, 32'd594, 32'd2919},
{-32'd1001, -32'd4294, 32'd3366, 32'd4374},
{-32'd6638, 32'd3065, -32'd374, 32'd5098},
{-32'd3933, 32'd3503, -32'd8455, 32'd2094},
{32'd2290, 32'd3591, 32'd718, 32'd6728},
{-32'd623, 32'd175, -32'd8417, -32'd902},
{32'd4015, -32'd87, 32'd4016, 32'd8043},
{32'd5390, -32'd628, 32'd5168, 32'd977},
{32'd3863, 32'd3643, 32'd1341, 32'd3407},
{-32'd406, -32'd8691, -32'd6495, -32'd1347},
{32'd5312, 32'd4809, -32'd582, 32'd6871},
{-32'd2427, 32'd4420, 32'd5114, -32'd2347},
{-32'd13058, -32'd8107, 32'd3316, -32'd3986},
{32'd11602, 32'd6073, 32'd3675, 32'd4896},
{-32'd5248, -32'd12357, -32'd7200, -32'd2469},
{-32'd10370, 32'd6281, -32'd9631, 32'd692},
{-32'd9900, -32'd1089, 32'd12045, -32'd2165},
{-32'd4927, 32'd8847, -32'd32, 32'd5940},
{-32'd9199, -32'd1671, 32'd806, -32'd262},
{32'd2569, -32'd11183, -32'd10148, -32'd176},
{32'd1928, -32'd2606, -32'd14, -32'd3371},
{32'd301, -32'd3094, 32'd36, -32'd5579},
{32'd9865, 32'd2725, -32'd1704, -32'd2954},
{-32'd1147, -32'd5991, -32'd3067, -32'd7440},
{-32'd1383, -32'd7352, 32'd4724, -32'd3061},
{-32'd1941, 32'd177, 32'd6599, 32'd5124},
{-32'd4281, 32'd6276, 32'd1415, -32'd796},
{-32'd3047, -32'd957, 32'd5142, 32'd2642},
{32'd2361, -32'd4877, 32'd691, -32'd5877},
{-32'd5026, 32'd404, -32'd7659, -32'd2540},
{32'd1771, 32'd7975, 32'd1131, 32'd2303},
{-32'd3816, -32'd4174, -32'd1574, -32'd2139},
{32'd10036, -32'd2388, 32'd2574, -32'd1615},
{32'd8188, 32'd7715, 32'd2196, -32'd3331},
{-32'd5886, 32'd3359, 32'd6089, -32'd1334},
{32'd186, 32'd410, 32'd3329, 32'd4506},
{-32'd1182, -32'd3990, -32'd742, -32'd6004},
{-32'd2544, -32'd2005, 32'd359, -32'd1406},
{32'd5181, 32'd654, 32'd1763, 32'd6260},
{32'd6585, 32'd4548, 32'd5445, 32'd2057},
{32'd2141, 32'd3312, -32'd7628, 32'd922},
{-32'd5460, -32'd6780, -32'd3227, -32'd3168},
{-32'd2413, -32'd5039, -32'd7812, 32'd3944},
{-32'd2982, 32'd5006, 32'd3902, -32'd3019},
{32'd2474, -32'd1238, 32'd5617, 32'd3283},
{-32'd3092, 32'd2490, 32'd2504, -32'd1190},
{-32'd8772, 32'd754, -32'd7350, 32'd871},
{32'd3795, -32'd558, 32'd6129, -32'd1693},
{-32'd1414, -32'd3453, 32'd1674, -32'd1798},
{32'd3474, 32'd3248, -32'd8708, -32'd1944},
{32'd1829, -32'd10713, 32'd3396, -32'd7415},
{-32'd4986, 32'd320, -32'd2218, -32'd4114},
{32'd519, 32'd44, 32'd807, 32'd4262},
{-32'd10667, -32'd2584, -32'd2580, -32'd1796},
{32'd5156, -32'd8329, 32'd2820, 32'd796},
{32'd5556, 32'd5118, 32'd2487, -32'd3192},
{32'd3942, 32'd1880, -32'd2130, -32'd1960},
{-32'd2512, 32'd4499, -32'd4984, 32'd2804},
{32'd2699, 32'd11391, 32'd6662, 32'd3174},
{32'd4142, 32'd1858, 32'd6618, -32'd5145},
{-32'd9083, -32'd395, -32'd6354, -32'd5899},
{32'd3436, -32'd6000, 32'd2186, -32'd6273},
{-32'd4000, 32'd13935, -32'd2611, 32'd3040},
{-32'd3644, 32'd14142, -32'd2181, -32'd1529},
{-32'd4053, 32'd2444, -32'd3880, -32'd6289},
{32'd5450, 32'd4971, 32'd522, -32'd224},
{32'd3718, -32'd4746, -32'd7446, -32'd1790},
{32'd1394, 32'd5959, 32'd4517, 32'd2383},
{-32'd13527, -32'd6974, -32'd5370, -32'd263},
{-32'd2430, -32'd7951, -32'd185, -32'd1675},
{32'd543, 32'd2294, 32'd1422, -32'd1426},
{-32'd1231, 32'd6375, -32'd1722, 32'd3209},
{-32'd2849, -32'd2067, -32'd6233, 32'd2996},
{32'd3078, 32'd501, 32'd3122, -32'd3046},
{32'd1171, -32'd7260, 32'd1528, 32'd1536},
{32'd7482, 32'd567, 32'd13178, -32'd5851},
{-32'd305, 32'd7635, -32'd1541, -32'd3535},
{32'd4504, 32'd1535, 32'd5959, 32'd2300},
{-32'd9504, 32'd1578, 32'd3947, 32'd2495},
{-32'd4634, -32'd6260, -32'd3928, 32'd148},
{32'd13172, -32'd4918, 32'd1922, 32'd2861},
{32'd5035, 32'd7225, -32'd2211, -32'd534},
{-32'd4389, 32'd7733, 32'd3514, -32'd408},
{-32'd844, -32'd5437, -32'd4877, 32'd593},
{-32'd4528, -32'd10726, -32'd40, 32'd2194},
{32'd3988, -32'd4732, -32'd1273, 32'd3056},
{32'd978, -32'd1792, 32'd1873, 32'd3358},
{32'd2063, -32'd4114, -32'd4412, -32'd1105},
{32'd998, 32'd9291, 32'd1384, -32'd3542},
{-32'd2743, -32'd2619, 32'd2596, -32'd531},
{-32'd1452, -32'd575, 32'd337, 32'd3464},
{-32'd3960, -32'd2189, -32'd1703, 32'd1440},
{-32'd4560, -32'd10283, 32'd3648, 32'd3209},
{-32'd4901, -32'd1006, -32'd5984, 32'd17},
{32'd6313, -32'd239, 32'd2058, 32'd782},
{-32'd3136, -32'd1642, -32'd4906, -32'd1953},
{-32'd158, -32'd202, -32'd2398, -32'd7001},
{-32'd1188, 32'd2813, -32'd5998, 32'd2542},
{-32'd745, 32'd2457, -32'd5785, -32'd653},
{32'd4352, 32'd4173, -32'd1724, 32'd7005},
{-32'd1444, 32'd558, 32'd4825, -32'd4852},
{32'd145, -32'd2466, -32'd2687, 32'd3380},
{-32'd129, -32'd10722, -32'd1838, -32'd214},
{32'd10342, 32'd6182, 32'd1723, -32'd7191},
{-32'd8440, 32'd6315, -32'd3451, -32'd957},
{-32'd5884, -32'd9666, -32'd1463, -32'd6158},
{32'd576, -32'd2518, -32'd4018, 32'd303},
{-32'd3748, -32'd3946, 32'd4135, 32'd379},
{-32'd2857, -32'd11089, -32'd3224, -32'd2255},
{-32'd1100, 32'd2016, 32'd4671, -32'd2371},
{32'd11, -32'd1565, -32'd154, -32'd5167},
{32'd3722, -32'd3687, -32'd3284, -32'd7425},
{-32'd1121, 32'd6762, -32'd2813, -32'd1852},
{32'd7149, -32'd6877, 32'd4148, -32'd333},
{-32'd9397, -32'd9757, -32'd3785, -32'd5712},
{32'd5465, -32'd4657, 32'd7006, -32'd113},
{32'd2572, 32'd1617, 32'd3948, 32'd3078},
{32'd4799, -32'd3899, 32'd3490, 32'd396},
{-32'd1483, -32'd1290, -32'd3412, -32'd290},
{-32'd2980, -32'd2053, 32'd3240, -32'd1653},
{32'd3467, -32'd4139, 32'd1470, 32'd2544},
{-32'd9329, 32'd2030, -32'd8255, 32'd2186},
{-32'd1663, 32'd2301, 32'd8050, 32'd1399},
{32'd4825, 32'd9287, 32'd9190, 32'd4268},
{-32'd1246, 32'd5529, -32'd5525, 32'd2936},
{32'd3097, 32'd3942, -32'd4532, -32'd508},
{-32'd243, -32'd7657, 32'd6829, -32'd4542},
{-32'd948, -32'd4210, 32'd3209, 32'd7778},
{32'd6238, 32'd5470, 32'd2736, -32'd3508},
{-32'd3301, 32'd1476, -32'd1355, -32'd3068},
{-32'd1696, -32'd5818, 32'd1970, -32'd5620},
{32'd5089, -32'd3646, -32'd7371, 32'd3458},
{-32'd10202, 32'd261, -32'd1863, -32'd4491},
{-32'd3708, -32'd3901, 32'd1928, 32'd1476},
{32'd1162, -32'd2891, -32'd824, 32'd381},
{32'd5105, 32'd1369, -32'd903, -32'd330},
{32'd2628, 32'd9603, -32'd10, 32'd2301},
{32'd5303, 32'd2253, -32'd2134, 32'd2678},
{32'd14198, -32'd6069, 32'd812, -32'd37},
{-32'd147, 32'd3222, 32'd2411, 32'd4322},
{32'd4973, -32'd1284, -32'd823, 32'd3496},
{-32'd5746, -32'd1682, -32'd2428, -32'd3743},
{-32'd1237, -32'd9489, -32'd5070, 32'd157},
{-32'd3953, 32'd793, 32'd6286, 32'd4168},
{-32'd4282, -32'd3106, 32'd2455, 32'd1360},
{32'd938, -32'd3837, 32'd1012, -32'd4705},
{32'd3602, 32'd3469, -32'd805, 32'd1155},
{32'd12246, -32'd6209, 32'd5472, -32'd2539},
{-32'd6473, -32'd7917, -32'd1962, -32'd4354},
{-32'd2660, -32'd9281, 32'd3218, -32'd4667},
{-32'd7684, -32'd961, -32'd1417, -32'd650},
{-32'd6725, 32'd2860, -32'd6871, -32'd2694},
{32'd6318, 32'd5480, -32'd3261, 32'd1817},
{-32'd2689, 32'd69, 32'd3760, 32'd1257},
{-32'd8266, -32'd126, 32'd627, -32'd3152},
{-32'd2995, 32'd2323, 32'd697, 32'd5640},
{-32'd2064, -32'd3085, -32'd5616, -32'd5379},
{-32'd2610, -32'd5528, -32'd5383, -32'd2755},
{32'd15207, 32'd2798, 32'd3148, 32'd4458},
{-32'd1780, 32'd8663, 32'd503, 32'd2415},
{32'd1260, -32'd93, -32'd494, -32'd115},
{32'd2505, 32'd7804, -32'd2362, 32'd6570},
{32'd11701, -32'd2157, -32'd192, 32'd6695},
{32'd3361, 32'd2982, -32'd2717, 32'd4464},
{-32'd4163, 32'd5411, -32'd3107, -32'd5229},
{32'd1408, -32'd2309, 32'd2525, 32'd814},
{-32'd696, 32'd7613, -32'd2423, 32'd965},
{-32'd210, -32'd2540, -32'd1189, 32'd4612},
{-32'd15, -32'd4133, -32'd2209, 32'd1303},
{32'd1783, -32'd2654, 32'd2712, 32'd2202},
{32'd5738, -32'd8327, -32'd4587, 32'd7223},
{-32'd3683, -32'd5301, 32'd418, -32'd565},
{-32'd3805, -32'd9139, -32'd8019, 32'd5867},
{-32'd388, 32'd1134, 32'd4550, -32'd2729},
{-32'd2959, -32'd13305, 32'd5705, 32'd5108},
{32'd8027, 32'd10435, 32'd2629, 32'd245},
{-32'd2641, 32'd7307, -32'd4493, 32'd2317},
{32'd2907, -32'd2525, -32'd535, -32'd1353},
{-32'd2154, -32'd4350, 32'd528, -32'd788},
{32'd5500, -32'd2269, 32'd2809, -32'd1685},
{32'd6945, -32'd2148, -32'd5115, 32'd3020},
{32'd2257, 32'd6142, 32'd5421, -32'd1133},
{-32'd14240, 32'd9478, -32'd271, 32'd4738},
{32'd5122, -32'd727, -32'd7129, -32'd2818},
{32'd3813, 32'd70, -32'd6157, 32'd6666},
{-32'd7313, -32'd2233, 32'd343, 32'd6081},
{-32'd6475, 32'd2411, 32'd7723, -32'd2105},
{32'd5052, -32'd2421, -32'd6612, -32'd6088},
{32'd8021, 32'd6458, -32'd6335, 32'd4474},
{32'd2115, 32'd6614, 32'd3039, 32'd426},
{32'd15302, 32'd6169, 32'd5532, 32'd6312},
{-32'd4095, -32'd3386, -32'd2560, 32'd2478},
{-32'd4992, 32'd1027, -32'd6880, -32'd3187},
{-32'd6773, -32'd2279, -32'd4692, -32'd5043},
{32'd2640, -32'd2042, 32'd9226, -32'd1872},
{32'd13706, -32'd2037, -32'd2871, 32'd1630},
{32'd12273, -32'd4671, -32'd2934, -32'd1480},
{-32'd7597, -32'd12745, 32'd26, 32'd2889},
{32'd2163, 32'd9202, 32'd1036, 32'd1397},
{-32'd4993, 32'd930, -32'd4591, -32'd586},
{32'd1682, -32'd889, -32'd279, 32'd3526},
{-32'd1805, 32'd1425, -32'd3605, -32'd6105},
{-32'd6171, 32'd1524, -32'd2331, -32'd2499},
{-32'd3392, -32'd3110, 32'd3533, 32'd4016},
{-32'd2982, -32'd3226, -32'd5869, -32'd934},
{32'd6193, -32'd1603, -32'd1993, 32'd3740},
{-32'd1809, -32'd3869, 32'd2754, -32'd4472},
{-32'd9914, 32'd2127, 32'd2824, -32'd3576},
{-32'd2856, -32'd7260, -32'd10913, -32'd6191},
{-32'd1551, 32'd4014, -32'd5266, -32'd5914},
{32'd7218, -32'd2116, 32'd2828, 32'd2363},
{32'd4148, 32'd330, 32'd4147, -32'd2273},
{-32'd3415, 32'd1663, 32'd1062, 32'd2104},
{32'd2090, 32'd187, 32'd4562, 32'd4005}
},
{{-32'd15710, -32'd7880, -32'd1207, -32'd879},
{32'd15256, -32'd2589, -32'd7433, 32'd5559},
{32'd6476, 32'd983, -32'd1451, 32'd7595},
{32'd20574, 32'd5182, 32'd7798, -32'd6712},
{32'd4691, 32'd19053, 32'd21299, 32'd1822},
{32'd651, -32'd3237, -32'd1881, -32'd1445},
{32'd9738, 32'd6657, 32'd20654, 32'd2375},
{-32'd2449, 32'd8162, 32'd793, -32'd2813},
{32'd18226, 32'd2546, 32'd371, -32'd2624},
{32'd6790, -32'd2362, 32'd15926, 32'd882},
{-32'd1394, -32'd2357, -32'd7163, 32'd3933},
{32'd3754, -32'd10557, 32'd481, 32'd125},
{-32'd12593, -32'd8285, 32'd3178, -32'd4799},
{32'd2333, 32'd3197, -32'd10181, 32'd6734},
{32'd2981, 32'd9538, -32'd16350, 32'd245},
{-32'd12009, -32'd3840, 32'd1400, -32'd16723},
{32'd3191, 32'd21105, 32'd1159, 32'd631},
{-32'd11081, -32'd10188, 32'd7308, 32'd18454},
{-32'd4512, 32'd2518, 32'd6308, -32'd8254},
{32'd2420, 32'd2227, 32'd6031, -32'd7525},
{-32'd7901, -32'd4618, 32'd4295, -32'd12274},
{-32'd408, -32'd2262, -32'd10739, -32'd5188},
{-32'd9748, 32'd1694, 32'd4487, 32'd175},
{32'd5956, -32'd2174, -32'd414, 32'd2692},
{-32'd10254, -32'd1320, 32'd15383, 32'd4884},
{-32'd8, 32'd1205, 32'd1428, -32'd1623},
{-32'd7928, -32'd7708, 32'd6067, -32'd11843},
{-32'd2497, 32'd3059, 32'd10762, -32'd1763},
{-32'd7092, -32'd15840, -32'd4411, -32'd13881},
{32'd8484, 32'd4956, 32'd2727, 32'd14479},
{-32'd10030, 32'd8398, -32'd522, -32'd10193},
{32'd1104, 32'd2423, -32'd3019, 32'd792},
{-32'd4867, 32'd9538, 32'd1226, 32'd364},
{-32'd5271, 32'd1182, 32'd2965, 32'd2366},
{32'd424, -32'd66, 32'd14968, 32'd6930},
{32'd6669, -32'd2076, -32'd2855, 32'd7400},
{-32'd672, -32'd3215, -32'd2116, -32'd4474},
{-32'd1205, 32'd10561, -32'd3761, -32'd11495},
{-32'd17627, -32'd4038, -32'd2365, -32'd1309},
{-32'd3386, 32'd346, -32'd509, 32'd10421},
{32'd1059, -32'd3774, -32'd10824, -32'd12772},
{32'd5528, -32'd241, 32'd3397, 32'd9908},
{-32'd3773, 32'd6154, 32'd7855, 32'd14119},
{-32'd1440, 32'd4670, -32'd2616, 32'd1271},
{-32'd7954, 32'd3444, -32'd7958, -32'd12366},
{-32'd14826, 32'd2540, 32'd1512, -32'd6390},
{-32'd1779, -32'd544, -32'd19884, -32'd16082},
{32'd108, -32'd579, -32'd10301, 32'd998},
{-32'd3741, -32'd12648, 32'd6421, 32'd2288},
{-32'd11338, 32'd754, -32'd13658, 32'd11443},
{32'd6694, -32'd44, 32'd2192, 32'd8705},
{32'd1456, 32'd1320, 32'd9442, 32'd3003},
{-32'd3729, 32'd351, -32'd898, -32'd11393},
{-32'd1201, 32'd3205, -32'd6742, 32'd13365},
{-32'd5786, 32'd13385, 32'd8913, -32'd1137},
{-32'd19750, 32'd471, -32'd17545, -32'd7475},
{-32'd13422, 32'd9419, -32'd2293, 32'd766},
{-32'd6297, -32'd838, -32'd9128, -32'd6676},
{32'd3822, -32'd8162, -32'd8456, -32'd352},
{-32'd13709, -32'd13443, 32'd6039, -32'd8002},
{-32'd2242, 32'd17692, -32'd712, -32'd1632},
{-32'd12700, 32'd6908, -32'd1933, 32'd7899},
{-32'd3465, -32'd7356, -32'd16092, -32'd3435},
{-32'd5810, -32'd7210, -32'd3670, -32'd6101},
{-32'd869, 32'd4749, -32'd10714, -32'd12606},
{-32'd182, -32'd3164, 32'd13830, 32'd9127},
{-32'd9748, 32'd7650, -32'd13232, -32'd19574},
{32'd13030, -32'd717, -32'd5405, 32'd1060},
{-32'd17208, -32'd7248, -32'd15573, -32'd14776},
{32'd5381, 32'd2267, 32'd7415, 32'd3550},
{32'd1111, -32'd8178, 32'd7645, -32'd8565},
{32'd8331, -32'd4196, 32'd2552, 32'd4418},
{-32'd14015, -32'd14578, -32'd4618, 32'd3953},
{32'd2443, 32'd11951, -32'd13284, 32'd2460},
{-32'd4236, 32'd1431, 32'd3538, 32'd8066},
{32'd2903, 32'd5967, 32'd4500, 32'd5401},
{32'd6477, 32'd13132, -32'd18003, 32'd320},
{-32'd584, 32'd1123, -32'd7, 32'd5741},
{32'd5646, 32'd9208, -32'd4847, -32'd4162},
{-32'd10831, 32'd5776, -32'd10305, 32'd3226},
{-32'd2572, 32'd3294, 32'd12798, -32'd1988},
{32'd5072, 32'd12060, 32'd9100, 32'd3837},
{-32'd14391, -32'd7291, -32'd17818, -32'd6918},
{32'd2249, 32'd6630, 32'd7736, 32'd10905},
{32'd1358, 32'd4685, 32'd37, 32'd10564},
{32'd3137, 32'd787, -32'd3254, -32'd12844},
{-32'd3416, 32'd5922, 32'd5422, 32'd14668},
{-32'd10811, -32'd5499, -32'd6069, -32'd147},
{-32'd7625, -32'd4069, 32'd4751, -32'd11993},
{-32'd1053, -32'd8886, 32'd609, -32'd14713},
{32'd4039, -32'd9597, 32'd9379, 32'd9556},
{-32'd2425, 32'd3744, 32'd1824, -32'd3063},
{32'd6861, 32'd1652, 32'd8599, 32'd4154},
{32'd3790, 32'd1599, 32'd10665, 32'd2866},
{-32'd3780, 32'd5899, 32'd979, -32'd11132},
{-32'd2528, -32'd1658, -32'd8717, -32'd4078},
{32'd10620, 32'd11156, 32'd11992, -32'd4421},
{-32'd1098, -32'd6936, 32'd15383, 32'd16196},
{32'd5224, 32'd10583, 32'd14559, 32'd2818},
{-32'd157, -32'd5003, 32'd8265, 32'd1889},
{32'd2846, -32'd13711, -32'd14471, -32'd5539},
{32'd8576, 32'd602, 32'd9946, 32'd3736},
{32'd2263, 32'd4277, -32'd11363, -32'd3856},
{-32'd5061, -32'd10235, 32'd7696, -32'd8110},
{-32'd27766, -32'd4767, -32'd7716, 32'd9975},
{32'd7266, 32'd696, 32'd5223, -32'd510},
{-32'd25952, 32'd5484, -32'd2280, 32'd2226},
{32'd9112, 32'd3915, -32'd5796, -32'd10077},
{32'd2020, -32'd11301, 32'd8895, -32'd6717},
{-32'd7869, -32'd325, -32'd130, 32'd4112},
{-32'd10490, 32'd15158, -32'd4679, -32'd1564},
{32'd402, -32'd7064, 32'd201, 32'd4496},
{-32'd9480, 32'd3894, -32'd1922, 32'd13936},
{-32'd9847, 32'd1918, 32'd3174, 32'd3367},
{-32'd3407, -32'd9262, -32'd9131, -32'd7029},
{-32'd3344, 32'd1273, -32'd3078, 32'd8205},
{32'd15936, -32'd9155, 32'd8990, 32'd8285},
{32'd30418, 32'd891, 32'd124, 32'd9609},
{32'd10476, 32'd25916, -32'd7314, -32'd1162},
{32'd11518, -32'd3325, 32'd7830, -32'd3600},
{-32'd4614, -32'd18363, 32'd5561, -32'd9419},
{32'd16167, 32'd9658, -32'd731, -32'd4189},
{32'd2626, -32'd4843, 32'd3059, -32'd240},
{32'd18473, -32'd368, 32'd8361, -32'd2130},
{-32'd17369, -32'd2450, 32'd11534, 32'd1393},
{-32'd8177, 32'd6005, 32'd4349, 32'd11483},
{32'd11388, -32'd20039, -32'd5576, -32'd10516},
{32'd1743, -32'd1454, -32'd12402, 32'd1746},
{-32'd2191, -32'd4936, -32'd29, -32'd14592},
{32'd331, -32'd4519, 32'd3244, -32'd410},
{-32'd1127, 32'd2216, -32'd3429, -32'd5133},
{32'd2661, -32'd472, -32'd2938, 32'd7984},
{-32'd10639, 32'd7297, -32'd8471, -32'd13736},
{32'd13600, 32'd2902, 32'd8134, 32'd2214},
{-32'd3032, -32'd8362, 32'd1546, -32'd5655},
{32'd3324, 32'd85, 32'd1928, -32'd1198},
{-32'd12680, 32'd6551, -32'd10353, 32'd9825},
{-32'd628, -32'd14481, -32'd405, 32'd1614},
{32'd7116, -32'd11571, 32'd6074, -32'd2735},
{-32'd8287, -32'd7393, -32'd16227, -32'd8885},
{32'd3060, -32'd3850, 32'd1264, 32'd17423},
{-32'd2382, -32'd250, 32'd6630, -32'd2790},
{32'd8943, -32'd4906, -32'd2735, 32'd13},
{32'd2425, 32'd6987, -32'd1170, -32'd10219},
{32'd15922, 32'd2172, 32'd5899, 32'd4011},
{32'd16654, 32'd10837, 32'd8347, 32'd15114},
{-32'd2521, 32'd2892, -32'd2511, 32'd5619},
{-32'd9457, 32'd8602, -32'd20961, -32'd11911},
{32'd17087, 32'd11913, 32'd12361, -32'd1857},
{-32'd13164, -32'd13119, -32'd9745, -32'd12923},
{-32'd10047, 32'd6575, -32'd12176, -32'd3590},
{-32'd3183, 32'd11309, 32'd4362, 32'd4917},
{-32'd11739, -32'd8067, 32'd2524, -32'd8451},
{32'd7564, -32'd660, -32'd11516, 32'd660},
{-32'd10109, 32'd1774, -32'd12573, 32'd5106},
{32'd19850, 32'd14959, 32'd1499, 32'd8826},
{-32'd16330, -32'd4774, 32'd1244, 32'd4791},
{-32'd13702, 32'd9391, -32'd1326, 32'd5305},
{32'd4259, 32'd1134, 32'd7493, -32'd17033},
{-32'd10029, -32'd15715, -32'd6611, -32'd2238},
{32'd11639, 32'd4241, -32'd2930, 32'd6186},
{-32'd1823, 32'd7497, 32'd1138, 32'd8259},
{32'd545, -32'd1829, -32'd14023, -32'd5489},
{32'd13887, 32'd6869, 32'd5574, 32'd17377},
{32'd1139, -32'd234, 32'd6109, -32'd4928},
{-32'd19385, -32'd3008, -32'd14981, -32'd6593},
{32'd4102, 32'd1814, 32'd5112, -32'd7845},
{-32'd795, 32'd5736, -32'd8761, -32'd16857},
{32'd4377, -32'd1615, -32'd2122, -32'd4984},
{-32'd776, 32'd9358, -32'd12691, -32'd7122},
{32'd2319, 32'd4128, -32'd2884, 32'd6673},
{32'd1116, 32'd3094, -32'd7437, -32'd4791},
{32'd1356, 32'd1282, 32'd12467, 32'd7162},
{32'd6197, 32'd8985, 32'd1195, -32'd10985},
{32'd9628, 32'd8576, 32'd9633, 32'd2363},
{-32'd20941, 32'd12844, -32'd1308, 32'd274},
{32'd6560, -32'd538, 32'd8656, 32'd19252},
{-32'd8679, -32'd11884, 32'd3204, -32'd11780},
{32'd2920, -32'd9351, 32'd3684, 32'd7524},
{-32'd9986, 32'd3496, -32'd15026, -32'd9772},
{32'd12257, 32'd5828, 32'd2770, -32'd2395},
{-32'd3057, -32'd2843, -32'd15656, -32'd3546},
{-32'd6167, 32'd3544, -32'd5225, -32'd2416},
{-32'd608, 32'd6107, 32'd7933, -32'd10144},
{-32'd697, 32'd1133, 32'd4026, -32'd1367},
{-32'd1107, -32'd7193, 32'd7039, -32'd12212},
{32'd16534, -32'd5460, 32'd1421, 32'd10278},
{32'd3666, 32'd11344, -32'd7243, 32'd7853},
{-32'd3956, 32'd3410, 32'd2773, 32'd10168},
{32'd2011, -32'd3422, -32'd9287, -32'd248},
{-32'd556, 32'd10832, 32'd7472, -32'd9254},
{32'd1380, -32'd4482, 32'd1719, 32'd10418},
{-32'd13996, -32'd12631, 32'd4574, -32'd3897},
{-32'd3841, -32'd3249, -32'd790, 32'd1537},
{32'd4343, -32'd18321, 32'd4031, -32'd8848},
{-32'd4456, -32'd8261, -32'd1161, -32'd4653},
{32'd2347, 32'd4268, -32'd12878, -32'd1608},
{32'd3461, 32'd2016, 32'd9469, -32'd9715},
{-32'd8769, 32'd139, -32'd13589, 32'd884},
{32'd13812, -32'd845, 32'd4658, -32'd1312},
{-32'd6367, -32'd3088, -32'd24127, -32'd2044},
{32'd481, 32'd6901, 32'd2354, -32'd10620},
{32'd2575, 32'd3683, 32'd10722, 32'd2890},
{-32'd2194, 32'd22253, 32'd1159, 32'd10417},
{-32'd20382, 32'd3242, -32'd5215, -32'd10830},
{32'd7903, -32'd8210, -32'd4407, -32'd678},
{-32'd4986, 32'd8151, -32'd1999, 32'd7704},
{32'd10566, -32'd2731, -32'd2760, -32'd11698},
{-32'd17116, 32'd6896, -32'd7434, 32'd1019},
{32'd1418, -32'd9564, 32'd9436, -32'd152},
{-32'd538, 32'd57, -32'd5433, 32'd441},
{-32'd24888, -32'd2237, 32'd12877, -32'd9489},
{32'd854, 32'd4823, -32'd5625, -32'd3016},
{-32'd5828, -32'd3687, 32'd1167, 32'd455},
{-32'd11624, 32'd1969, 32'd3144, -32'd7323},
{-32'd8296, 32'd6187, 32'd7946, 32'd3159},
{32'd7895, 32'd7898, -32'd1575, 32'd5038},
{32'd4017, 32'd5514, 32'd3530, -32'd12825},
{32'd8048, 32'd1851, 32'd1667, -32'd2117},
{32'd7343, 32'd11385, 32'd1528, -32'd5407},
{-32'd3408, 32'd5485, -32'd4904, 32'd11287},
{-32'd7291, -32'd5588, 32'd520, 32'd706},
{-32'd6992, -32'd12257, 32'd13162, 32'd2838},
{32'd1997, -32'd14342, -32'd12274, -32'd6327},
{-32'd20915, -32'd7805, 32'd6116, -32'd9120},
{-32'd984, 32'd2745, -32'd2849, 32'd10352},
{32'd6394, 32'd1499, -32'd1783, 32'd3539},
{32'd2351, -32'd9036, 32'd6840, 32'd1883},
{-32'd5997, 32'd1561, 32'd10640, -32'd2492},
{32'd2775, 32'd1220, 32'd1626, -32'd164},
{32'd5671, -32'd14739, -32'd5425, 32'd5747},
{32'd9567, 32'd897, 32'd5021, 32'd1506},
{-32'd285, -32'd4078, 32'd3751, -32'd7396},
{32'd5258, -32'd5979, 32'd2255, 32'd12669},
{-32'd718, 32'd7742, 32'd2724, -32'd2711},
{-32'd1527, 32'd3201, -32'd10962, 32'd7623},
{32'd3633, -32'd5035, 32'd4261, -32'd2625},
{32'd3774, 32'd6176, -32'd3452, 32'd2701},
{32'd3397, 32'd4561, 32'd4877, -32'd1270},
{32'd2978, -32'd6710, 32'd8242, -32'd15754},
{32'd11109, -32'd9086, -32'd10470, -32'd18},
{32'd3724, 32'd12814, 32'd5865, -32'd1143},
{-32'd5307, 32'd1645, -32'd8071, 32'd397},
{32'd4571, 32'd11198, 32'd4276, 32'd1828},
{-32'd3667, -32'd2086, 32'd9176, 32'd2006},
{-32'd24, 32'd8257, -32'd16853, 32'd5897},
{32'd2757, 32'd6490, -32'd10293, -32'd6967},
{-32'd12074, -32'd11107, 32'd520, -32'd7846},
{32'd3485, 32'd1272, -32'd2002, 32'd11915},
{-32'd13275, 32'd12859, -32'd2521, -32'd8957},
{32'd9186, 32'd12079, -32'd2590, -32'd5805},
{-32'd1667, 32'd3285, -32'd5750, 32'd5847},
{32'd7121, 32'd6058, 32'd6803, -32'd2809},
{-32'd7363, 32'd5870, -32'd5525, -32'd3766},
{-32'd2774, 32'd3966, -32'd9198, 32'd7379},
{32'd13630, -32'd1112, 32'd306, 32'd8799},
{32'd5027, -32'd2041, -32'd4971, -32'd7743},
{32'd4189, 32'd347, 32'd11619, -32'd1121},
{32'd6345, -32'd2728, -32'd4843, -32'd236},
{-32'd527, 32'd5600, 32'd5063, 32'd3048},
{32'd16605, -32'd3064, 32'd3455, 32'd1023},
{-32'd2295, -32'd6959, 32'd3062, -32'd8612},
{32'd3254, 32'd18759, -32'd3314, -32'd2312},
{-32'd1390, -32'd5143, -32'd807, 32'd2263},
{32'd3894, 32'd784, 32'd9138, 32'd11879},
{32'd6240, -32'd9813, -32'd186, 32'd6854},
{32'd14995, -32'd8499, 32'd3282, 32'd699},
{-32'd10778, -32'd1682, -32'd9372, -32'd700},
{32'd443, 32'd2945, -32'd7212, 32'd1789},
{32'd2093, 32'd5642, -32'd18504, -32'd7093},
{-32'd16806, -32'd5686, 32'd3216, 32'd100},
{-32'd7018, 32'd2269, 32'd15192, 32'd13332},
{-32'd19143, -32'd246, -32'd12769, 32'd873},
{-32'd6711, 32'd13145, -32'd1236, 32'd8800},
{32'd13013, 32'd15568, 32'd4592, -32'd4872},
{-32'd18025, -32'd8144, -32'd6925, 32'd4846},
{32'd8089, -32'd573, 32'd21669, 32'd4913},
{32'd10112, -32'd5921, 32'd6613, -32'd13747},
{-32'd6592, 32'd3841, 32'd41, 32'd942},
{32'd7014, -32'd513, -32'd1325, -32'd2879},
{-32'd7377, 32'd3423, 32'd1343, -32'd4222},
{-32'd5052, 32'd6634, -32'd4359, 32'd8245},
{32'd704, 32'd3136, -32'd2785, -32'd12163},
{32'd878, 32'd5348, 32'd5627, -32'd157},
{32'd752, -32'd6675, 32'd11389, 32'd11693},
{-32'd13942, 32'd10333, -32'd14204, -32'd4382},
{-32'd4301, -32'd1463, 32'd5005, -32'd2561},
{32'd6007, 32'd1155, -32'd3708, -32'd3967},
{32'd3837, 32'd6722, 32'd8537, 32'd2471},
{32'd9566, -32'd11031, -32'd10452, 32'd21652},
{32'd8046, -32'd6373, 32'd5023, 32'd7487},
{-32'd5176, -32'd2825, 32'd13369, -32'd2774},
{-32'd5614, -32'd18189, -32'd8495, 32'd3212},
{-32'd9444, -32'd12808, -32'd577, 32'd11634},
{32'd959, -32'd17381, -32'd8464, 32'd3557},
{-32'd10255, 32'd4181, -32'd5743, 32'd5517},
{32'd10777, 32'd754, -32'd3740, 32'd3753},
{32'd308, 32'd312, 32'd3321, -32'd5466},
{32'd7829, 32'd4962, 32'd7500, -32'd1023},
{-32'd17498, -32'd16039, 32'd403, -32'd4217}
},
{{32'd7492, 32'd6532, 32'd7295, 32'd3861},
{-32'd356, 32'd3425, -32'd3060, -32'd10032},
{32'd4366, 32'd3691, -32'd6007, 32'd4200},
{32'd11352, -32'd150, 32'd2883, 32'd4456},
{32'd1363, 32'd9334, 32'd6150, -32'd820},
{32'd1592, 32'd718, 32'd6112, 32'd484},
{-32'd5088, 32'd6749, -32'd3303, 32'd12782},
{-32'd7040, -32'd4300, -32'd1926, -32'd16630},
{-32'd10814, -32'd7262, -32'd9921, -32'd3464},
{32'd10698, 32'd9375, 32'd5125, 32'd5977},
{-32'd5181, 32'd3981, 32'd2048, 32'd1083},
{32'd2183, -32'd1187, -32'd5271, -32'd3444},
{32'd8578, -32'd314, -32'd12606, 32'd1270},
{32'd4374, -32'd4501, -32'd3872, 32'd3216},
{32'd1565, -32'd4629, -32'd4574, 32'd9846},
{32'd2031, -32'd2353, -32'd774, -32'd5806},
{32'd7551, -32'd1347, 32'd2217, -32'd662},
{32'd4249, 32'd3789, 32'd5538, -32'd1705},
{32'd5194, 32'd5267, 32'd2826, -32'd5256},
{-32'd3599, 32'd2453, -32'd3504, -32'd3827},
{32'd3235, 32'd2224, -32'd6727, -32'd3126},
{-32'd3314, -32'd5658, -32'd11640, -32'd7445},
{-32'd2033, -32'd4392, -32'd11921, -32'd15699},
{32'd6587, -32'd6502, -32'd783, 32'd1369},
{32'd3834, 32'd6514, 32'd4726, 32'd3062},
{32'd555, -32'd9134, -32'd5926, -32'd1625},
{-32'd6167, -32'd3854, 32'd1794, 32'd168},
{-32'd8332, 32'd1974, -32'd2181, -32'd3496},
{32'd6898, 32'd814, 32'd8425, -32'd6491},
{-32'd4232, -32'd923, 32'd695, 32'd3477},
{32'd111, -32'd3983, -32'd11757, -32'd9448},
{-32'd9222, -32'd933, -32'd949, 32'd5655},
{-32'd2579, 32'd5392, 32'd10464, -32'd6749},
{32'd1313, -32'd8328, -32'd3010, -32'd4225},
{32'd5960, 32'd5722, 32'd6749, 32'd7259},
{32'd3477, -32'd2560, 32'd3718, 32'd4065},
{-32'd4382, -32'd2228, 32'd5883, -32'd5322},
{32'd6999, -32'd3668, 32'd46, 32'd1353},
{32'd4535, -32'd1793, 32'd102, 32'd1051},
{-32'd3496, 32'd2040, 32'd5932, 32'd6244},
{-32'd269, 32'd4417, -32'd1260, 32'd3560},
{32'd2901, 32'd8596, 32'd4960, 32'd5929},
{32'd5252, -32'd912, -32'd1616, 32'd109},
{-32'd5316, -32'd4413, -32'd8030, -32'd6652},
{-32'd5993, -32'd7412, -32'd9687, -32'd12330},
{-32'd4434, 32'd2106, 32'd915, -32'd4327},
{-32'd1275, 32'd802, -32'd3917, -32'd8507},
{-32'd3482, -32'd2956, 32'd8797, -32'd840},
{-32'd302, -32'd4422, 32'd8603, -32'd1864},
{-32'd3485, 32'd5191, -32'd10469, -32'd5301},
{-32'd6067, 32'd2769, -32'd11465, -32'd7136},
{32'd4763, -32'd3761, 32'd8418, 32'd12051},
{-32'd2199, -32'd2402, 32'd659, 32'd4147},
{-32'd3438, -32'd921, -32'd2378, 32'd4635},
{-32'd2813, -32'd3975, -32'd3213, -32'd2067},
{-32'd780, -32'd3910, -32'd3283, -32'd7936},
{32'd6032, 32'd5452, 32'd11920, 32'd7940},
{-32'd22482, -32'd3013, -32'd1376, -32'd7456},
{-32'd5583, -32'd4349, -32'd4368, -32'd854},
{-32'd5501, -32'd3957, 32'd6191, -32'd552},
{-32'd7566, -32'd4249, 32'd3308, -32'd533},
{-32'd18415, 32'd3156, 32'd12389, 32'd10419},
{-32'd7008, -32'd2380, -32'd1645, 32'd2975},
{-32'd7867, -32'd6385, 32'd785, 32'd8370},
{-32'd447, -32'd3164, 32'd5, -32'd4379},
{32'd874, 32'd1225, 32'd7839, 32'd6144},
{-32'd7054, -32'd922, -32'd3266, 32'd3919},
{-32'd4249, -32'd2229, 32'd6247, -32'd7653},
{-32'd3160, 32'd6792, -32'd3993, -32'd10793},
{-32'd6739, 32'd896, 32'd9260, 32'd5069},
{-32'd4978, -32'd1374, -32'd2444, -32'd6006},
{32'd7357, 32'd4457, -32'd103, 32'd3652},
{-32'd8166, 32'd5580, -32'd6439, -32'd4380},
{32'd4008, -32'd107, -32'd2825, -32'd3861},
{-32'd5987, -32'd2210, 32'd6796, 32'd2119},
{-32'd2359, 32'd381, -32'd3566, 32'd6480},
{-32'd6181, 32'd2639, -32'd18352, -32'd6300},
{-32'd2278, -32'd14385, -32'd3559, 32'd2991},
{32'd1236, 32'd5159, -32'd2585, -32'd860},
{32'd5749, 32'd1818, 32'd13162, 32'd3677},
{-32'd3381, 32'd4721, 32'd1380, -32'd4151},
{-32'd2013, 32'd5200, 32'd6584, 32'd2286},
{-32'd501, 32'd2394, 32'd7631, -32'd7579},
{32'd1983, 32'd5073, -32'd2257, 32'd7242},
{32'd731, -32'd500, -32'd8516, -32'd2334},
{-32'd6954, -32'd2806, 32'd11935, -32'd3101},
{32'd8255, -32'd6672, 32'd4205, 32'd9273},
{-32'd2516, -32'd12001, -32'd8852, -32'd10369},
{-32'd5587, -32'd1061, -32'd7380, -32'd5282},
{32'd403, -32'd4063, 32'd2475, -32'd1775},
{32'd1144, 32'd6584, 32'd5939, -32'd1556},
{-32'd4744, 32'd3052, 32'd0, -32'd1530},
{-32'd25, 32'd7472, 32'd569, -32'd8498},
{32'd6143, 32'd159, 32'd4013, 32'd2263},
{-32'd2988, -32'd556, 32'd5534, 32'd85},
{-32'd3652, 32'd8015, -32'd2510, -32'd1306},
{32'd10693, 32'd6917, 32'd6604, 32'd2947},
{-32'd2558, 32'd2373, 32'd469, 32'd7070},
{32'd9119, 32'd1291, 32'd3420, 32'd3100},
{32'd6674, 32'd8992, 32'd6134, -32'd2017},
{-32'd8153, -32'd4551, -32'd6963, 32'd816},
{-32'd4399, 32'd3643, -32'd11698, -32'd3591},
{-32'd3891, 32'd7797, 32'd2558, 32'd3421},
{-32'd386, -32'd5772, 32'd1373, 32'd7936},
{32'd772, 32'd3863, 32'd5067, 32'd11531},
{-32'd5197, -32'd4051, 32'd2419, 32'd2819},
{-32'd7217, 32'd2340, -32'd3245, 32'd797},
{32'd2052, -32'd5399, -32'd7214, 32'd1836},
{32'd8427, 32'd6538, -32'd2271, -32'd1717},
{32'd3415, 32'd64, -32'd7581, -32'd3123},
{-32'd5400, 32'd5593, -32'd4715, -32'd1819},
{-32'd2640, 32'd2713, 32'd7009, -32'd975},
{-32'd1448, 32'd828, -32'd2959, -32'd2526},
{-32'd1807, 32'd4569, 32'd5159, 32'd3245},
{32'd2426, 32'd604, 32'd2490, -32'd947},
{-32'd10149, 32'd1216, -32'd4746, 32'd147},
{32'd9452, 32'd4678, -32'd3919, -32'd934},
{32'd1949, 32'd4301, -32'd1092, -32'd2074},
{32'd89, 32'd5349, 32'd1235, -32'd4813},
{32'd120, 32'd6174, 32'd17827, 32'd16799},
{32'd2297, -32'd3281, 32'd3726, -32'd897},
{-32'd7794, 32'd5992, -32'd1501, 32'd9914},
{-32'd1278, 32'd3199, 32'd5567, -32'd1239},
{32'd1158, 32'd7533, -32'd1684, 32'd537},
{-32'd6703, -32'd5410, -32'd1740, -32'd5144},
{-32'd2399, -32'd577, -32'd9289, -32'd603},
{-32'd8016, 32'd2499, -32'd2267, -32'd839},
{-32'd5029, -32'd1080, -32'd576, -32'd11975},
{32'd4214, -32'd2425, -32'd3290, -32'd6105},
{-32'd5900, -32'd5585, -32'd2796, -32'd781},
{32'd1259, 32'd3143, 32'd5488, 32'd7145},
{32'd2623, -32'd810, -32'd10590, -32'd7685},
{-32'd21999, -32'd3894, -32'd12315, -32'd3869},
{-32'd1670, 32'd3099, 32'd5464, 32'd1129},
{32'd7500, 32'd7674, 32'd868, -32'd9950},
{-32'd1364, 32'd6178, 32'd706, -32'd6156},
{-32'd6261, 32'd416, 32'd1131, -32'd8015},
{32'd5140, -32'd4703, -32'd9392, -32'd4494},
{-32'd6698, -32'd4881, 32'd4577, -32'd2235},
{-32'd9775, -32'd13553, 32'd859, 32'd944},
{32'd8897, 32'd6706, 32'd2266, 32'd8960},
{32'd5074, -32'd3013, -32'd2031, -32'd2141},
{32'd514, 32'd883, 32'd6759, -32'd215},
{-32'd7348, -32'd830, -32'd5619, -32'd3298},
{-32'd554, 32'd6477, 32'd5119, 32'd13621},
{32'd4899, 32'd2192, -32'd3085, -32'd2112},
{-32'd46, -32'd3613, -32'd11435, -32'd8596},
{32'd3991, 32'd7537, 32'd1356, 32'd2125},
{-32'd254, -32'd3552, 32'd3649, 32'd10291},
{32'd6963, -32'd1285, 32'd8879, -32'd4553},
{-32'd3852, -32'd5154, -32'd7672, -32'd4236},
{32'd7822, 32'd2990, -32'd1670, -32'd2096},
{-32'd6470, -32'd6402, 32'd8499, -32'd472},
{32'd7375, -32'd1741, -32'd4, 32'd1023},
{32'd187, -32'd2515, -32'd7312, -32'd9629},
{-32'd4644, -32'd6056, 32'd921, 32'd6398},
{32'd8079, 32'd6677, -32'd9050, -32'd6318},
{32'd5977, -32'd342, 32'd5763, 32'd3103},
{-32'd8041, -32'd8343, -32'd558, 32'd279},
{32'd9632, 32'd10523, 32'd1467, 32'd406},
{32'd4982, -32'd4723, 32'd3127, 32'd6214},
{-32'd3113, 32'd4162, 32'd4098, -32'd740},
{-32'd6559, -32'd480, -32'd6496, 32'd704},
{-32'd2140, 32'd6126, -32'd2856, 32'd11347},
{-32'd717, 32'd1230, 32'd51, -32'd583},
{-32'd3259, 32'd5966, 32'd3451, 32'd2543},
{-32'd1636, -32'd540, -32'd2079, 32'd1492},
{32'd508, -32'd2785, -32'd6992, -32'd11545},
{32'd1729, -32'd2979, 32'd5659, 32'd4081},
{-32'd10521, -32'd14343, 32'd8050, 32'd7421},
{32'd4571, -32'd4218, -32'd2300, 32'd12882},
{-32'd1142, -32'd1471, 32'd8938, 32'd1074},
{32'd9355, 32'd6341, 32'd4889, 32'd2006},
{-32'd10590, -32'd83, -32'd2774, 32'd9787},
{32'd6708, 32'd2839, -32'd5509, 32'd1178},
{32'd849, -32'd1928, 32'd6255, -32'd605},
{-32'd679, 32'd3441, 32'd968, -32'd2254},
{-32'd3892, -32'd2242, -32'd9597, -32'd6264},
{32'd4877, 32'd2205, 32'd1373, -32'd3302},
{-32'd1477, -32'd3130, -32'd7209, -32'd6099},
{-32'd6384, 32'd2497, -32'd8082, 32'd2310},
{-32'd662, -32'd1750, 32'd4012, 32'd26},
{-32'd223, -32'd1871, 32'd1672, -32'd3232},
{-32'd4702, -32'd4251, 32'd573, 32'd3153},
{32'd4210, -32'd4323, -32'd1705, -32'd9129},
{-32'd21, 32'd4776, 32'd6697, -32'd31},
{32'd1210, 32'd8337, 32'd242, 32'd9761},
{32'd5530, -32'd2936, 32'd3993, -32'd1855},
{-32'd4069, -32'd6249, -32'd1707, -32'd3100},
{-32'd3171, 32'd11639, -32'd8285, -32'd8713},
{32'd882, 32'd5182, 32'd8568, 32'd638},
{32'd3939, -32'd4486, -32'd4624, 32'd6716},
{-32'd2325, -32'd7660, 32'd5764, 32'd1312},
{32'd408, -32'd3340, 32'd3213, -32'd10253},
{32'd5891, -32'd7778, -32'd4216, -32'd2748},
{32'd1570, -32'd721, 32'd1534, -32'd2614},
{32'd1671, 32'd3775, -32'd4353, -32'd5885},
{32'd10757, -32'd2238, 32'd1861, -32'd2032},
{32'd695, 32'd6057, -32'd7397, -32'd7622},
{-32'd6563, 32'd1217, -32'd829, -32'd4129},
{-32'd7327, -32'd3268, -32'd6674, -32'd5104},
{-32'd7955, 32'd461, 32'd5829, -32'd3617},
{-32'd658, 32'd1466, 32'd6833, -32'd274},
{32'd6901, 32'd819, -32'd466, 32'd7129},
{-32'd7773, -32'd7072, -32'd8076, -32'd5102},
{32'd6240, 32'd3448, 32'd1615, 32'd507},
{32'd2103, 32'd1161, -32'd101, 32'd3351},
{-32'd3243, -32'd5369, -32'd8263, -32'd3091},
{32'd808, -32'd1058, -32'd2213, 32'd3938},
{-32'd324, 32'd4056, 32'd1358, 32'd5350},
{-32'd4861, -32'd1828, 32'd5795, -32'd1983},
{32'd1707, -32'd5947, -32'd1725, 32'd5239},
{32'd1282, -32'd2008, -32'd4817, -32'd8447},
{32'd2233, 32'd5244, 32'd7070, 32'd2551},
{32'd3409, -32'd4492, -32'd16968, 32'd468},
{32'd1619, 32'd138, 32'd8212, 32'd7466},
{32'd5905, -32'd8443, 32'd697, -32'd1182},
{32'd4166, -32'd6320, -32'd18440, -32'd8303},
{-32'd969, 32'd886, 32'd9085, 32'd12247},
{-32'd6936, -32'd3833, -32'd5831, -32'd3899},
{-32'd3261, -32'd4837, -32'd12713, -32'd6826},
{-32'd2265, 32'd4714, -32'd4742, 32'd5374},
{-32'd3327, 32'd621, 32'd4800, -32'd751},
{-32'd3054, -32'd2440, 32'd4010, -32'd2340},
{32'd5377, 32'd5512, 32'd6015, -32'd2754},
{-32'd1855, -32'd2414, 32'd7778, 32'd8565},
{32'd2247, 32'd321, -32'd5998, -32'd16722},
{-32'd5077, -32'd2126, -32'd2785, -32'd5732},
{32'd4375, 32'd3040, 32'd334, -32'd4308},
{32'd8184, 32'd5822, 32'd8594, 32'd61},
{-32'd2484, 32'd98, 32'd3437, -32'd71},
{-32'd10371, -32'd115, 32'd915, 32'd2325},
{32'd3288, 32'd2340, 32'd4316, 32'd6698},
{-32'd1597, 32'd4661, -32'd6482, 32'd2585},
{-32'd3588, -32'd1510, -32'd2584, -32'd9917},
{-32'd2458, 32'd2010, -32'd1642, -32'd8019},
{32'd8680, 32'd3251, 32'd11209, -32'd2749},
{-32'd5879, 32'd1930, -32'd10527, -32'd565},
{32'd6371, 32'd2297, 32'd444, -32'd5223},
{-32'd9709, -32'd1281, -32'd1977, 32'd905},
{32'd6303, -32'd442, 32'd5844, -32'd4068},
{-32'd4733, -32'd2577, -32'd9361, -32'd934},
{-32'd3032, -32'd7292, -32'd8767, -32'd6278},
{32'd7552, -32'd5302, -32'd11117, 32'd3395},
{32'd3897, 32'd8058, 32'd5394, -32'd3054},
{32'd1619, 32'd5241, 32'd3770, 32'd3753},
{32'd595, -32'd1825, -32'd6206, 32'd5296},
{-32'd3405, 32'd2901, 32'd6629, -32'd4238},
{-32'd395, -32'd2260, 32'd6310, 32'd897},
{32'd7831, -32'd5147, 32'd1005, 32'd5423},
{-32'd8812, -32'd9637, -32'd3446, -32'd3535},
{-32'd210, 32'd8365, 32'd1508, 32'd1592},
{32'd727, 32'd683, -32'd617, -32'd6770},
{32'd1472, -32'd4221, -32'd2106, -32'd1286},
{-32'd3750, -32'd3057, -32'd3029, 32'd15},
{32'd2779, 32'd145, 32'd12808, 32'd6900},
{32'd1554, 32'd1524, 32'd10195, -32'd4114},
{32'd4444, 32'd2637, 32'd3468, 32'd5665},
{-32'd5584, -32'd5298, -32'd3937, 32'd4676},
{-32'd1128, -32'd3011, 32'd6497, 32'd1174},
{-32'd2782, -32'd2325, 32'd5570, 32'd2844},
{32'd3327, 32'd1869, -32'd2, -32'd1142},
{-32'd499, 32'd1471, -32'd1579, -32'd418},
{32'd3487, -32'd2542, -32'd7151, 32'd236},
{-32'd3944, -32'd2355, 32'd982, 32'd421},
{-32'd8989, 32'd3183, 32'd7954, 32'd5001},
{32'd8296, 32'd10828, 32'd2159, 32'd2998},
{-32'd3107, 32'd1692, -32'd1638, -32'd10314},
{32'd809, 32'd2282, 32'd304, -32'd3871},
{32'd189, -32'd1690, -32'd1766, 32'd7430},
{32'd11548, -32'd2794, 32'd1746, -32'd5918},
{32'd5129, -32'd1570, 32'd1284, 32'd3166},
{-32'd11524, 32'd1909, 32'd14416, 32'd1947},
{-32'd6691, -32'd4414, -32'd2924, -32'd747},
{32'd12410, -32'd3503, -32'd3839, -32'd6735},
{-32'd2081, 32'd3484, -32'd9516, -32'd4345},
{32'd10835, 32'd8781, 32'd6461, 32'd7111},
{32'd6096, -32'd1595, -32'd1546, 32'd118},
{-32'd5657, -32'd9431, -32'd6363, -32'd6808},
{-32'd1317, -32'd3756, -32'd6496, -32'd387},
{-32'd5569, -32'd1075, 32'd8621, -32'd3038},
{-32'd3775, 32'd1942, -32'd14296, -32'd3381},
{32'd3885, 32'd2403, -32'd5899, -32'd2935},
{-32'd1118, -32'd290, 32'd669, 32'd10481},
{32'd1784, -32'd6538, 32'd2778, -32'd4556},
{-32'd5535, -32'd4407, -32'd15103, -32'd3628},
{32'd38, 32'd5478, -32'd1669, -32'd1390},
{-32'd1679, -32'd4270, -32'd999, 32'd3046},
{32'd6934, 32'd4427, -32'd5069, 32'd9442},
{-32'd7780, 32'd12922, 32'd2451, 32'd2159},
{-32'd9064, 32'd2229, -32'd4148, -32'd2588},
{32'd7187, 32'd9995, 32'd9080, 32'd7319},
{-32'd1546, -32'd3127, -32'd10860, 32'd163},
{-32'd2299, -32'd4104, -32'd7596, 32'd2149},
{32'd2686, -32'd2538, -32'd5730, 32'd489},
{32'd887, -32'd4970, -32'd5627, -32'd798},
{-32'd8483, -32'd484, -32'd5823, 32'd7012},
{32'd8628, -32'd550, 32'd4521, 32'd4461},
{32'd9806, 32'd2572, -32'd3924, 32'd7583},
{32'd3507, 32'd706, -32'd865, -32'd6013}
},
{{-32'd298, 32'd6081, 32'd7106, 32'd1637},
{-32'd6371, -32'd2442, -32'd5147, -32'd6121},
{-32'd8709, 32'd4583, 32'd5441, -32'd5037},
{-32'd2784, 32'd249, 32'd3024, 32'd4257},
{32'd7749, 32'd78, 32'd7485, 32'd7051},
{32'd8062, 32'd6710, 32'd1290, -32'd1184},
{32'd3537, 32'd7340, 32'd2967, -32'd11380},
{-32'd12917, -32'd2342, -32'd611, -32'd8272},
{-32'd8318, 32'd1363, -32'd9525, 32'd842},
{32'd8349, 32'd15106, -32'd1795, 32'd4474},
{-32'd6702, -32'd4043, 32'd3397, -32'd140},
{-32'd8651, -32'd2569, -32'd5388, 32'd7151},
{32'd1635, 32'd12663, 32'd6555, -32'd4883},
{32'd5149, 32'd3596, -32'd5482, 32'd5282},
{-32'd15066, 32'd2393, -32'd7728, 32'd291},
{-32'd3365, 32'd3245, 32'd2402, -32'd4705},
{-32'd284, -32'd3676, 32'd3342, 32'd6260},
{-32'd3391, 32'd89, 32'd3786, -32'd2163},
{32'd3063, 32'd19089, -32'd182, -32'd352},
{32'd7661, -32'd5491, -32'd11831, 32'd2808},
{32'd6182, 32'd4103, -32'd5126, 32'd214},
{32'd1556, -32'd9751, 32'd4455, 32'd317},
{32'd2748, -32'd12759, -32'd4616, -32'd4702},
{-32'd2923, -32'd1831, -32'd5433, -32'd13261},
{32'd865, 32'd16963, 32'd3142, 32'd8089},
{32'd2628, 32'd12508, -32'd7009, -32'd4907},
{32'd12160, 32'd4136, -32'd4372, 32'd8746},
{-32'd2641, 32'd4261, -32'd3542, -32'd14836},
{-32'd10068, 32'd9472, 32'd13157, 32'd9783},
{-32'd10887, 32'd4343, -32'd2395, 32'd14033},
{32'd158, 32'd11228, -32'd6707, 32'd15668},
{-32'd2136, 32'd7488, -32'd9335, -32'd2082},
{32'd1191, 32'd14771, 32'd9845, -32'd81},
{32'd538, 32'd2355, 32'd8617, 32'd2060},
{32'd6187, 32'd11716, -32'd3511, -32'd379},
{-32'd4153, -32'd4590, -32'd7833, 32'd5487},
{-32'd1966, 32'd8181, -32'd12772, 32'd120},
{-32'd7292, -32'd1712, 32'd382, -32'd17330},
{-32'd4000, 32'd3214, -32'd484, -32'd1847},
{-32'd5969, -32'd5170, 32'd6673, -32'd2926},
{-32'd1948, -32'd1695, -32'd3909, 32'd3985},
{32'd8679, 32'd8486, -32'd76, -32'd599},
{-32'd73, -32'd1094, -32'd2108, -32'd15860},
{32'd2589, 32'd184, -32'd3609, -32'd13673},
{32'd684, -32'd10104, -32'd4988, -32'd8581},
{-32'd1149, -32'd3171, -32'd2824, 32'd9523},
{-32'd13819, -32'd191, -32'd5949, -32'd4988},
{-32'd8523, -32'd2755, -32'd3017, 32'd6594},
{32'd223, 32'd3515, 32'd10169, -32'd2305},
{-32'd342, 32'd5895, -32'd1727, -32'd9125},
{32'd9321, -32'd4914, 32'd5014, 32'd13114},
{32'd640, 32'd8658, 32'd7678, -32'd5710},
{32'd1880, 32'd2963, -32'd14459, -32'd3889},
{-32'd2072, -32'd9290, -32'd10695, -32'd6645},
{-32'd253, 32'd7662, 32'd1593, -32'd714},
{32'd1225, -32'd5199, -32'd5559, 32'd5641},
{-32'd12907, 32'd16226, -32'd1812, 32'd7162},
{-32'd2757, 32'd6220, 32'd4132, -32'd5830},
{-32'd3813, -32'd7327, -32'd1485, -32'd4987},
{-32'd1063, -32'd4411, -32'd16333, 32'd9035},
{32'd10400, -32'd8295, -32'd4743, 32'd11872},
{-32'd5331, -32'd3732, 32'd7898, 32'd4285},
{-32'd4585, -32'd17612, -32'd3582, -32'd129},
{32'd9657, 32'd5490, -32'd14388, 32'd4015},
{-32'd6222, -32'd6065, -32'd4613, -32'd8706},
{-32'd71, 32'd11063, -32'd6466, -32'd962},
{-32'd331, 32'd6103, -32'd9241, 32'd8938},
{-32'd7245, -32'd10785, -32'd13411, -32'd11149},
{-32'd5523, -32'd3936, 32'd8108, 32'd4012},
{-32'd3991, -32'd4485, 32'd6019, 32'd4948},
{-32'd4725, -32'd724, -32'd3636, 32'd3193},
{-32'd1605, 32'd6675, 32'd6495, -32'd5388},
{-32'd801, -32'd3053, -32'd6890, 32'd2083},
{32'd4681, -32'd5685, 32'd13732, 32'd4617},
{32'd10125, 32'd5932, 32'd12468, -32'd1008},
{-32'd1522, -32'd12509, -32'd3900, -32'd7604},
{-32'd7085, 32'd2708, 32'd4161, -32'd4804},
{32'd3723, -32'd7741, 32'd11423, 32'd12262},
{-32'd775, 32'd8849, -32'd6790, 32'd66},
{32'd2199, -32'd6446, 32'd12797, 32'd5109},
{-32'd4618, 32'd6651, -32'd5679, 32'd565},
{32'd6218, -32'd15179, -32'd3809, -32'd2658},
{-32'd7431, 32'd4806, 32'd6509, 32'd5582},
{32'd11904, -32'd6021, 32'd3197, 32'd3469},
{-32'd6453, -32'd3840, 32'd4051, -32'd4770},
{-32'd10637, -32'd8202, -32'd12908, 32'd9976},
{32'd1173, -32'd8834, -32'd5196, -32'd5968},
{32'd409, -32'd10141, -32'd185, 32'd3392},
{-32'd1544, -32'd2703, 32'd5108, 32'd9348},
{-32'd5847, -32'd7953, -32'd6449, 32'd10065},
{32'd5340, 32'd4814, -32'd3295, -32'd2321},
{-32'd1829, -32'd3140, -32'd2020, 32'd3667},
{-32'd2676, 32'd8637, -32'd5294, -32'd7151},
{32'd1842, 32'd6528, 32'd2589, -32'd4060},
{-32'd8051, -32'd3632, 32'd859, -32'd632},
{-32'd4488, -32'd9052, -32'd4849, -32'd7218},
{32'd3806, 32'd12956, -32'd4003, -32'd2615},
{32'd1538, 32'd3234, 32'd10369, -32'd6966},
{-32'd1785, 32'd2439, -32'd3063, -32'd3085},
{32'd6105, 32'd7587, 32'd6591, 32'd5072},
{-32'd11830, -32'd1344, -32'd19292, -32'd13596},
{-32'd6558, -32'd2982, -32'd12028, 32'd4103},
{-32'd3051, -32'd6788, -32'd58, -32'd13114},
{32'd883, -32'd7821, 32'd545, 32'd3643},
{32'd2692, 32'd2413, -32'd2081, -32'd7636},
{32'd2379, 32'd5010, 32'd1180, 32'd1580},
{32'd5932, 32'd1978, -32'd7424, -32'd2227},
{-32'd6950, 32'd3766, 32'd4091, 32'd850},
{-32'd6385, 32'd1192, -32'd9637, -32'd1341},
{-32'd7106, -32'd7838, -32'd10458, -32'd5457},
{-32'd1006, -32'd8652, -32'd2175, 32'd3325},
{-32'd1886, -32'd8826, 32'd2123, -32'd5903},
{32'd1774, -32'd2677, 32'd8914, 32'd3796},
{-32'd5586, 32'd96, 32'd1719, 32'd2472},
{-32'd5341, -32'd13431, 32'd5867, 32'd4673},
{32'd15357, -32'd3878, -32'd6777, 32'd2439},
{-32'd7295, -32'd6885, 32'd7741, 32'd432},
{-32'd5849, -32'd1632, -32'd3624, 32'd3754},
{32'd1438, 32'd7943, 32'd2606, 32'd3956},
{32'd10120, 32'd10102, -32'd996, 32'd3358},
{-32'd10688, -32'd1820, 32'd4838, 32'd3941},
{32'd9277, 32'd181, -32'd3038, -32'd3815},
{32'd2791, 32'd4727, 32'd7337, 32'd1370},
{-32'd600, -32'd8207, -32'd7438, 32'd98},
{-32'd4583, 32'd16966, 32'd5497, 32'd6703},
{32'd493, 32'd2395, -32'd1386, -32'd5051},
{32'd1356, -32'd2848, 32'd5663, -32'd6003},
{-32'd13333, -32'd6515, -32'd1986, 32'd4862},
{32'd7157, -32'd9019, -32'd5406, -32'd6087},
{32'd1589, -32'd2196, 32'd14543, -32'd7969},
{32'd824, -32'd1705, 32'd248, 32'd3375},
{-32'd2811, -32'd6247, 32'd589, -32'd6539},
{-32'd5714, -32'd9258, -32'd7016, -32'd4279},
{-32'd6179, 32'd5632, 32'd2897, 32'd158},
{-32'd6652, -32'd3276, 32'd4659, 32'd13509},
{-32'd5655, 32'd4837, -32'd343, 32'd3330},
{32'd1302, 32'd9913, -32'd1332, -32'd674},
{32'd8927, -32'd16075, -32'd7845, -32'd1804},
{-32'd8, 32'd9171, 32'd6714, -32'd734},
{32'd2229, -32'd14396, -32'd3611, -32'd15603},
{32'd22241, -32'd4816, 32'd7729, 32'd9707},
{32'd1887, 32'd2538, 32'd3161, 32'd116},
{32'd11814, -32'd1589, 32'd7346, 32'd1730},
{32'd79, 32'd10003, -32'd6692, -32'd10243},
{-32'd3826, -32'd1545, -32'd6995, 32'd2542},
{32'd14833, 32'd3763, 32'd13829, 32'd3163},
{-32'd205, -32'd8027, 32'd1641, -32'd12216},
{-32'd13593, 32'd9492, -32'd8888, 32'd7879},
{32'd7383, -32'd1155, -32'd1582, 32'd3186},
{-32'd13124, 32'd2753, 32'd2829, -32'd3520},
{-32'd7652, -32'd5750, 32'd5730, -32'd14125},
{32'd8108, 32'd1670, 32'd4321, 32'd997},
{-32'd6218, -32'd7751, -32'd5217, -32'd6578},
{32'd7445, -32'd127, 32'd14409, 32'd4623},
{-32'd16083, -32'd12677, -32'd3315, -32'd4513},
{32'd2380, 32'd10785, -32'd7042, -32'd7909},
{32'd5024, 32'd3906, -32'd1309, 32'd5468},
{-32'd14128, -32'd1776, 32'd10056, 32'd4441},
{-32'd10339, 32'd596, -32'd3780, -32'd8159},
{-32'd189, 32'd6121, 32'd2210, 32'd2169},
{-32'd8655, 32'd1562, -32'd335, 32'd12546},
{32'd1039, 32'd2065, -32'd2194, 32'd3479},
{32'd2059, -32'd8196, 32'd605, 32'd22},
{32'd6093, 32'd5061, 32'd12646, -32'd14},
{32'd8799, 32'd863, 32'd12298, -32'd7247},
{-32'd4158, 32'd2960, -32'd3086, 32'd2748},
{-32'd13151, 32'd1643, -32'd3579, -32'd5096},
{-32'd4077, 32'd2602, -32'd6620, 32'd2673},
{-32'd775, -32'd6868, -32'd3219, 32'd4008},
{-32'd12806, -32'd7304, 32'd10582, -32'd3124},
{-32'd4802, -32'd6744, 32'd2503, -32'd4327},
{32'd4410, 32'd11947, -32'd1685, -32'd12107},
{32'd6432, 32'd3203, -32'd7677, 32'd3184},
{-32'd15937, 32'd1410, -32'd2149, -32'd5599},
{-32'd576, 32'd4901, 32'd5096, 32'd813},
{32'd2514, -32'd6878, 32'd7937, 32'd4424},
{-32'd1734, -32'd3037, 32'd11711, 32'd8633},
{-32'd3201, 32'd9139, 32'd7573, -32'd1179},
{-32'd2361, 32'd567, 32'd4467, 32'd539},
{-32'd3903, -32'd5126, 32'd11608, -32'd9305},
{32'd94, -32'd12097, -32'd1326, 32'd12128},
{32'd877, -32'd5059, 32'd1855, -32'd5199},
{-32'd4900, -32'd3567, -32'd52, -32'd3281},
{-32'd2964, -32'd2371, 32'd14072, -32'd5846},
{-32'd16146, -32'd6570, -32'd430, -32'd8150},
{32'd5448, -32'd5505, 32'd1999, 32'd2918},
{32'd3404, 32'd9659, -32'd425, 32'd3982},
{32'd4470, 32'd6226, 32'd6295, -32'd4838},
{-32'd4086, 32'd3968, -32'd2573, 32'd546},
{32'd2360, 32'd7321, -32'd1499, -32'd384},
{32'd6892, 32'd3084, -32'd4328, -32'd11951},
{32'd3966, 32'd6109, -32'd6916, -32'd4330},
{-32'd5663, 32'd9733, -32'd11131, 32'd6233},
{-32'd3796, 32'd16996, -32'd10788, -32'd9052},
{-32'd5160, -32'd11867, -32'd8065, -32'd6028},
{32'd9612, 32'd2623, 32'd3395, 32'd3355},
{-32'd2137, -32'd12956, -32'd3253, -32'd11807},
{32'd10945, -32'd5848, 32'd8579, 32'd2863},
{32'd3341, 32'd2866, 32'd4433, -32'd388},
{-32'd30, 32'd3109, -32'd3090, 32'd1776},
{-32'd3881, -32'd12667, 32'd2131, -32'd4787},
{-32'd3635, 32'd2708, 32'd5928, 32'd4228},
{32'd5829, 32'd3787, 32'd17085, -32'd1456},
{32'd16130, 32'd8007, -32'd366, 32'd4902},
{-32'd2249, 32'd2244, -32'd3884, -32'd3790},
{-32'd8515, -32'd750, 32'd4220, -32'd9652},
{32'd19414, 32'd3421, -32'd562, -32'd273},
{-32'd1428, -32'd5667, 32'd4300, -32'd727},
{-32'd9404, 32'd709, 32'd82, 32'd3188},
{-32'd12052, -32'd1383, -32'd799, 32'd5629},
{-32'd1391, -32'd11388, -32'd6651, -32'd4821},
{-32'd382, -32'd8479, -32'd5522, 32'd6574},
{32'd4632, 32'd8655, -32'd1423, -32'd2417},
{32'd3279, -32'd2394, 32'd6024, -32'd11056},
{-32'd3868, 32'd4287, 32'd5007, 32'd903},
{-32'd183, 32'd6905, 32'd3502, 32'd4102},
{-32'd3564, -32'd12951, -32'd5198, -32'd6371},
{-32'd5769, -32'd228, -32'd1322, 32'd1959},
{-32'd3877, -32'd4357, 32'd7776, 32'd6162},
{-32'd11017, 32'd1691, 32'd8341, -32'd11071},
{32'd8196, -32'd7331, 32'd15480, -32'd141},
{32'd1239, -32'd42, -32'd1813, 32'd4463},
{32'd111, 32'd2220, -32'd2430, -32'd10146},
{32'd444, 32'd8227, 32'd13095, 32'd694},
{32'd1080, -32'd8096, -32'd5078, 32'd14614},
{32'd2395, -32'd18210, 32'd12186, -32'd6628},
{32'd461, 32'd1709, 32'd11356, -32'd389},
{-32'd3123, -32'd3000, -32'd4998, -32'd2674},
{32'd4287, -32'd439, 32'd9735, 32'd10744},
{-32'd2724, 32'd4410, -32'd13010, 32'd4505},
{-32'd2497, 32'd384, 32'd10694, 32'd8642},
{-32'd7208, -32'd5391, -32'd8426, 32'd2354},
{32'd9093, 32'd5362, 32'd15822, 32'd1839},
{-32'd5786, 32'd2929, -32'd10007, 32'd2205},
{-32'd239, -32'd94, 32'd7696, -32'd7843},
{-32'd7773, -32'd17911, -32'd6514, -32'd7479},
{-32'd8187, 32'd1819, -32'd3038, 32'd6410},
{32'd3346, -32'd2217, -32'd5978, -32'd8505},
{32'd1094, -32'd2908, 32'd9125, 32'd2816},
{-32'd1914, 32'd1978, -32'd162, -32'd6885},
{-32'd12983, -32'd328, -32'd7464, 32'd13136},
{32'd7396, -32'd6786, 32'd2718, -32'd1994},
{-32'd8073, -32'd12533, -32'd3986, -32'd3393},
{32'd1587, -32'd4912, -32'd6835, -32'd4493},
{32'd10051, 32'd14182, 32'd768, 32'd2666},
{32'd2978, 32'd6283, 32'd1123, 32'd10921},
{-32'd5443, 32'd1241, -32'd1320, -32'd20201},
{-32'd7064, 32'd3995, 32'd1453, 32'd6673},
{-32'd9807, -32'd3922, 32'd4249, -32'd1555},
{-32'd6078, -32'd11407, -32'd10018, -32'd1512},
{32'd2310, -32'd9895, -32'd55, -32'd7497},
{32'd8826, 32'd4375, -32'd3443, 32'd5951},
{32'd9016, 32'd3208, -32'd8147, 32'd3395},
{32'd1123, 32'd1727, 32'd4414, -32'd451},
{32'd7711, -32'd7764, 32'd10030, -32'd5934},
{-32'd3219, 32'd8609, -32'd2561, 32'd6067},
{32'd934, 32'd3765, -32'd6772, 32'd597},
{32'd9440, -32'd5100, 32'd6639, 32'd3737},
{-32'd14121, 32'd1907, 32'd3311, -32'd1292},
{32'd6348, -32'd8908, 32'd7845, -32'd1991},
{32'd775, 32'd1015, -32'd6061, -32'd1083},
{32'd1415, 32'd8063, -32'd2925, -32'd6581},
{32'd8957, -32'd11033, -32'd9342, -32'd2247},
{-32'd5415, -32'd3744, 32'd5971, 32'd4728},
{32'd3547, -32'd10600, 32'd12203, -32'd266},
{-32'd21526, -32'd5676, 32'd398, 32'd6437},
{32'd6579, 32'd10749, 32'd11952, 32'd5436},
{-32'd12851, 32'd6448, -32'd69, -32'd578},
{-32'd5099, -32'd1944, -32'd634, -32'd5930},
{32'd2626, -32'd1014, -32'd11427, -32'd3442},
{-32'd3032, -32'd9259, 32'd6829, 32'd10742},
{32'd1972, 32'd4787, -32'd1297, 32'd2443},
{-32'd7477, -32'd5541, -32'd1730, 32'd2045},
{32'd4515, -32'd9405, 32'd3102, 32'd7782},
{32'd832, -32'd8560, 32'd5821, 32'd12038},
{32'd7845, 32'd1744, -32'd6173, 32'd2754},
{32'd8902, 32'd16126, 32'd9, 32'd5893},
{-32'd6030, -32'd5945, -32'd4498, -32'd208},
{-32'd6899, -32'd10170, -32'd433, 32'd2900},
{-32'd10202, -32'd1303, -32'd7145, 32'd242},
{32'd5167, 32'd10270, -32'd6114, 32'd3145},
{-32'd415, -32'd4672, 32'd1529, -32'd7099},
{32'd10374, -32'd4516, 32'd5068, 32'd9256},
{32'd3989, 32'd2475, 32'd5148, 32'd5168},
{-32'd5912, -32'd2150, 32'd16055, 32'd6194},
{-32'd8207, -32'd11285, -32'd8264, -32'd10609},
{32'd8044, 32'd1592, -32'd6310, 32'd2941},
{32'd3035, -32'd10856, -32'd8876, -32'd10184},
{-32'd3104, -32'd6443, -32'd1794, -32'd5727},
{-32'd1951, -32'd2671, -32'd9236, -32'd3955},
{32'd8584, 32'd3184, 32'd6035, -32'd12563},
{32'd2205, 32'd10147, 32'd7352, 32'd5344},
{32'd5179, -32'd7241, -32'd3644, -32'd2913},
{32'd1917, -32'd1964, 32'd307, -32'd4288},
{-32'd6058, -32'd670, -32'd3691, 32'd8237},
{-32'd10266, -32'd8978, 32'd10277, -32'd4221},
{32'd4846, -32'd1657, 32'd5546, 32'd305},
{32'd5466, 32'd7941, -32'd4328, 32'd2731},
{32'd3312, 32'd16774, -32'd9580, 32'd6478},
{-32'd4181, 32'd9218, -32'd1214, 32'd6008}
},
{{32'd2908, 32'd3492, -32'd2000, 32'd5730},
{-32'd9848, -32'd4681, -32'd1407, 32'd2185},
{32'd9051, -32'd7716, -32'd8144, 32'd6151},
{-32'd8084, -32'd2024, 32'd6670, -32'd5586},
{32'd11808, 32'd1871, 32'd4457, 32'd2027},
{32'd248, -32'd5765, -32'd1128, 32'd4941},
{-32'd69, 32'd5340, 32'd11872, -32'd8533},
{-32'd3324, -32'd2684, -32'd3467, -32'd1856},
{-32'd9213, -32'd3728, 32'd3526, -32'd172},
{32'd13416, 32'd10820, 32'd8240, 32'd3131},
{-32'd1166, -32'd5851, 32'd3000, 32'd6571},
{32'd5122, 32'd9304, 32'd6446, 32'd3076},
{-32'd1180, 32'd4663, 32'd1683, -32'd4930},
{-32'd3030, -32'd6854, -32'd8442, -32'd7179},
{-32'd10853, -32'd3990, -32'd7584, -32'd9008},
{-32'd4125, -32'd12618, -32'd704, -32'd10558},
{32'd10530, -32'd9875, 32'd11083, -32'd5654},
{-32'd4095, 32'd2576, 32'd2808, -32'd2779},
{-32'd416, 32'd13007, -32'd4447, -32'd5983},
{-32'd3079, -32'd1578, 32'd6192, -32'd1391},
{-32'd1778, -32'd1249, -32'd1771, -32'd540},
{-32'd5903, -32'd3819, -32'd890, 32'd1607},
{-32'd6204, -32'd10384, -32'd3114, -32'd2636},
{-32'd11491, 32'd2789, -32'd6374, -32'd3379},
{32'd4989, 32'd10872, -32'd4562, 32'd8315},
{32'd3588, 32'd3845, -32'd6203, -32'd3428},
{-32'd816, -32'd9291, 32'd4085, 32'd15440},
{32'd4339, 32'd1719, -32'd4424, -32'd599},
{32'd126, 32'd12137, 32'd1421, -32'd1352},
{-32'd9540, 32'd9058, 32'd13657, -32'd1409},
{32'd35, -32'd10202, 32'd9146, 32'd5709},
{-32'd7813, -32'd13801, -32'd1950, 32'd6904},
{32'd15138, 32'd4499, -32'd7796, 32'd2302},
{32'd714, 32'd2475, -32'd11043, -32'd95},
{32'd10101, 32'd3949, 32'd10904, 32'd4421},
{32'd2413, -32'd13476, -32'd13106, 32'd5468},
{32'd5462, 32'd8321, -32'd1375, -32'd9071},
{-32'd7872, 32'd3936, -32'd489, -32'd7130},
{-32'd209, -32'd518, 32'd4553, 32'd5758},
{-32'd3520, 32'd2102, -32'd400, 32'd11273},
{32'd3162, -32'd277, 32'd3387, -32'd1571},
{32'd4073, -32'd732, -32'd1349, 32'd5208},
{-32'd8607, 32'd3573, 32'd4438, 32'd6303},
{-32'd3080, 32'd6167, -32'd4924, -32'd2579},
{32'd6665, 32'd2335, -32'd746, 32'd1448},
{32'd3184, -32'd862, 32'd78, 32'd2554},
{-32'd13039, -32'd3602, 32'd6887, -32'd6013},
{-32'd1475, -32'd9725, 32'd2392, 32'd1004},
{-32'd3182, 32'd1418, 32'd7611, -32'd4495},
{-32'd7119, -32'd2721, 32'd1477, -32'd4193},
{-32'd9159, -32'd8993, 32'd2235, 32'd6998},
{32'd3154, 32'd8076, 32'd2663, -32'd2950},
{-32'd660, -32'd14436, -32'd5101, -32'd3771},
{-32'd1029, 32'd5718, -32'd8614, -32'd3863},
{-32'd2498, 32'd11169, -32'd6255, -32'd2380},
{-32'd7794, -32'd7087, -32'd2101, -32'd66},
{32'd1486, 32'd5602, -32'd2252, 32'd10879},
{32'd2986, -32'd7513, 32'd2230, -32'd1728},
{-32'd1474, 32'd2042, 32'd12031, 32'd1718},
{32'd771, -32'd4181, 32'd1736, 32'd5006},
{-32'd976, -32'd6639, 32'd2031, 32'd7721},
{-32'd9603, 32'd1761, -32'd68, 32'd1106},
{-32'd6092, -32'd11732, 32'd605, -32'd2801},
{-32'd243, -32'd6047, -32'd1264, 32'd1108},
{32'd6764, 32'd10715, -32'd5881, -32'd7326},
{32'd11166, 32'd2364, 32'd3438, 32'd6659},
{-32'd6720, 32'd5650, 32'd12353, 32'd4007},
{-32'd3074, -32'd4438, 32'd5995, -32'd2610},
{-32'd4722, 32'd1696, -32'd8320, -32'd1628},
{32'd3000, 32'd6161, 32'd12990, -32'd1261},
{32'd11434, 32'd5365, -32'd2745, 32'd3066},
{-32'd287, 32'd5602, -32'd5668, -32'd989},
{-32'd9936, 32'd2326, -32'd6078, -32'd577},
{-32'd8351, -32'd921, 32'd8515, -32'd636},
{32'd5891, 32'd8906, -32'd3534, 32'd5217},
{-32'd585, 32'd398, 32'd1602, 32'd9585},
{32'd4370, -32'd4811, -32'd3171, -32'd5273},
{-32'd3024, 32'd1293, -32'd7948, -32'd99},
{32'd8760, 32'd2282, 32'd5608, -32'd3422},
{32'd1602, -32'd28, 32'd412, -32'd640},
{32'd11559, -32'd6833, 32'd4822, -32'd442},
{32'd13523, -32'd5707, 32'd1502, 32'd2456},
{-32'd2290, 32'd4735, -32'd1545, -32'd4864},
{32'd2979, 32'd261, 32'd10040, 32'd8573},
{-32'd2961, -32'd5998, -32'd2831, -32'd446},
{32'd4851, -32'd6145, 32'd2896, -32'd1521},
{32'd1711, 32'd10667, -32'd2627, -32'd2585},
{-32'd6238, -32'd4448, -32'd3860, -32'd12904},
{-32'd6098, -32'd4808, -32'd2031, 32'd3206},
{32'd479, -32'd3471, -32'd14104, -32'd1270},
{32'd105, 32'd8720, 32'd10622, -32'd994},
{-32'd10973, -32'd4090, -32'd132, 32'd1669},
{32'd3751, 32'd1037, -32'd3386, -32'd5927},
{32'd4727, -32'd10202, 32'd12803, -32'd8338},
{-32'd1917, -32'd3777, -32'd6574, -32'd4519},
{32'd4343, 32'd4650, -32'd231, -32'd731},
{32'd1932, 32'd8331, 32'd3045, -32'd6973},
{32'd781, -32'd3879, -32'd9563, 32'd4912},
{32'd7788, 32'd2826, 32'd3149, -32'd3716},
{32'd7855, 32'd145, 32'd9437, 32'd4899},
{32'd3394, -32'd5213, 32'd1688, -32'd7759},
{32'd1040, -32'd9597, 32'd13757, 32'd1626},
{32'd2017, 32'd7858, 32'd9432, -32'd8794},
{32'd9786, 32'd11718, 32'd5371, -32'd2130},
{-32'd348, 32'd4289, 32'd4775, 32'd1542},
{-32'd5894, -32'd8426, 32'd5798, 32'd3826},
{-32'd3881, -32'd4729, -32'd820, 32'd4574},
{-32'd3754, -32'd3689, -32'd5711, 32'd2335},
{32'd922, -32'd377, 32'd3249, 32'd402},
{-32'd6209, -32'd11487, -32'd3356, -32'd5544},
{32'd3308, 32'd8386, 32'd292, -32'd6727},
{32'd5496, 32'd11086, -32'd3601, -32'd4754},
{32'd10327, 32'd7338, -32'd6470, -32'd1523},
{32'd1506, -32'd5150, 32'd6974, 32'd8187},
{-32'd8241, -32'd9289, -32'd3952, 32'd3771},
{-32'd9470, -32'd6976, -32'd2075, 32'd343},
{32'd507, 32'd3777, 32'd11634, -32'd3442},
{32'd315, -32'd3343, -32'd168, -32'd3479},
{32'd5523, -32'd10344, 32'd8365, -32'd5825},
{32'd2990, -32'd106, 32'd161, 32'd7945},
{32'd3359, -32'd348, -32'd5614, 32'd10501},
{-32'd3799, 32'd10241, -32'd3367, -32'd230},
{32'd3259, -32'd5329, -32'd14146, 32'd6477},
{-32'd9244, -32'd2999, 32'd3439, 32'd1341},
{32'd839, 32'd3130, -32'd3962, 32'd15842},
{-32'd4443, 32'd8334, 32'd7543, -32'd637},
{-32'd3863, -32'd9216, 32'd5209, 32'd2359},
{32'd3924, -32'd5034, -32'd3276, 32'd4032},
{-32'd1110, 32'd3597, 32'd428, 32'd7167},
{32'd8400, 32'd617, -32'd7819, -32'd26},
{-32'd9783, -32'd1729, -32'd7900, -32'd1590},
{-32'd2002, 32'd6039, 32'd37, 32'd237},
{-32'd7887, -32'd5464, 32'd5937, -32'd7499},
{32'd2889, -32'd8128, 32'd6522, -32'd4602},
{32'd4119, 32'd8397, -32'd540, -32'd1101},
{32'd7829, -32'd8477, -32'd12495, -32'd445},
{32'd1636, 32'd3337, -32'd17361, 32'd1594},
{-32'd8830, 32'd3679, -32'd316, 32'd1609},
{32'd2596, -32'd985, -32'd2472, 32'd10146},
{-32'd2267, -32'd6438, -32'd3583, 32'd6244},
{32'd7846, 32'd3081, 32'd6582, -32'd3760},
{32'd8614, -32'd8129, -32'd12220, 32'd4864},
{32'd5217, 32'd2327, 32'd4641, 32'd4265},
{32'd2595, -32'd12344, 32'd3521, 32'd396},
{32'd5386, -32'd1123, -32'd1212, 32'd469},
{32'd6487, -32'd315, 32'd7578, 32'd564},
{-32'd2983, -32'd1080, -32'd950, 32'd2234},
{32'd2002, -32'd10671, 32'd303, 32'd9124},
{32'd9201, -32'd4488, 32'd4989, -32'd3774},
{-32'd9252, -32'd7127, -32'd5758, 32'd1247},
{-32'd6940, 32'd2997, -32'd9641, -32'd3020},
{32'd460, -32'd2937, 32'd5931, -32'd4599},
{32'd5883, -32'd3863, -32'd8117, 32'd4502},
{32'd6218, 32'd1231, 32'd1334, 32'd75},
{-32'd6194, 32'd6136, -32'd2577, 32'd283},
{32'd7968, -32'd2908, 32'd3607, -32'd1734},
{32'd683, 32'd1399, -32'd6748, 32'd5289},
{32'd778, 32'd3275, 32'd10303, -32'd4997},
{32'd2312, 32'd1388, 32'd1454, 32'd3335},
{-32'd7404, 32'd3219, -32'd15034, 32'd5706},
{-32'd16321, -32'd5344, -32'd2619, -32'd4966},
{32'd7031, -32'd930, -32'd4429, 32'd6409},
{-32'd5747, 32'd1593, 32'd1541, -32'd35},
{32'd14108, 32'd4583, 32'd19266, 32'd4314},
{32'd6777, 32'd1263, 32'd1952, 32'd3334},
{-32'd8399, -32'd1007, -32'd1900, 32'd4587},
{-32'd7958, -32'd1075, 32'd13877, -32'd3141},
{-32'd932, 32'd738, -32'd10910, 32'd13293},
{32'd1596, -32'd3834, -32'd432, -32'd11287},
{32'd2440, -32'd11681, -32'd1910, -32'd6240},
{-32'd6820, -32'd2888, 32'd566, 32'd4465},
{-32'd6307, 32'd5256, 32'd4429, 32'd619},
{32'd7381, 32'd8865, 32'd4897, -32'd4323},
{-32'd3046, -32'd7580, -32'd4811, -32'd12440},
{32'd6738, -32'd2446, 32'd1463, -32'd3100},
{32'd5179, 32'd7378, 32'd7638, 32'd2782},
{32'd7696, 32'd1131, 32'd7639, 32'd7076},
{-32'd2038, 32'd143, -32'd1574, 32'd2648},
{-32'd7551, -32'd5825, 32'd12617, 32'd3634},
{-32'd11834, -32'd8417, -32'd1834, 32'd6445},
{-32'd11718, -32'd6507, -32'd7297, 32'd2497},
{-32'd4713, -32'd5206, -32'd11554, 32'd1116},
{-32'd300, 32'd2241, 32'd692, 32'd1752},
{-32'd2474, -32'd2938, 32'd2057, 32'd4091},
{32'd3694, 32'd3475, 32'd2498, -32'd219},
{32'd8325, -32'd1227, 32'd7542, 32'd4877},
{32'd2340, 32'd1694, 32'd7835, 32'd4586},
{-32'd6544, -32'd2444, 32'd6440, -32'd239},
{32'd5437, -32'd8987, 32'd1373, -32'd6625},
{-32'd6747, 32'd5742, -32'd21113, 32'd744},
{-32'd6456, 32'd511, 32'd11013, -32'd3396},
{-32'd4723, -32'd2346, -32'd3780, -32'd1985},
{32'd1700, 32'd2707, 32'd2056, -32'd882},
{32'd2267, -32'd1638, 32'd4195, -32'd9020},
{-32'd987, 32'd2333, -32'd11304, -32'd3128},
{-32'd199, -32'd6050, -32'd8782, 32'd8287},
{-32'd541, -32'd887, 32'd1727, 32'd10723},
{32'd10280, 32'd11813, 32'd988, 32'd3886},
{32'd1832, 32'd515, 32'd393, 32'd3156},
{32'd5397, 32'd7886, 32'd11984, 32'd751},
{-32'd10287, -32'd4882, -32'd9314, -32'd4677},
{32'd949, 32'd1934, -32'd1357, -32'd4250},
{32'd5683, -32'd750, 32'd1672, 32'd7012},
{32'd4611, 32'd842, 32'd1649, -32'd1759},
{-32'd4216, -32'd3156, -32'd1165, 32'd1153},
{32'd757, 32'd7947, 32'd170, 32'd2281},
{32'd3763, -32'd9027, -32'd4144, 32'd4516},
{-32'd2025, -32'd3596, 32'd2833, -32'd3023},
{-32'd5007, -32'd6220, -32'd3811, 32'd5753},
{32'd9652, 32'd6499, 32'd3587, 32'd5176},
{32'd4032, 32'd4843, -32'd3282, -32'd5264},
{32'd3035, 32'd6733, 32'd990, 32'd3745},
{-32'd4005, -32'd9207, -32'd2028, 32'd5871},
{32'd4322, 32'd4431, 32'd950, -32'd3857},
{-32'd6047, 32'd940, -32'd5873, -32'd3127},
{-32'd8649, -32'd1726, -32'd274, -32'd5301},
{-32'd5693, -32'd9315, -32'd1960, -32'd7203},
{32'd4167, -32'd4343, -32'd332, 32'd6223},
{32'd1276, 32'd15053, -32'd1248, 32'd11441},
{-32'd8353, -32'd1779, 32'd6256, 32'd1114},
{-32'd10067, -32'd8827, 32'd3621, 32'd281},
{32'd679, 32'd79, 32'd9852, -32'd1116},
{32'd5588, 32'd1100, 32'd7552, 32'd1692},
{32'd8286, 32'd4932, -32'd2602, 32'd3490},
{32'd1568, -32'd4318, -32'd3551, 32'd8889},
{32'd2657, -32'd3649, -32'd2930, -32'd10614},
{-32'd6027, -32'd3529, -32'd7078, 32'd1491},
{32'd12563, -32'd5642, 32'd3098, -32'd882},
{32'd5078, -32'd5547, 32'd3489, -32'd6916},
{32'd6202, 32'd13142, 32'd719, -32'd3096},
{-32'd6756, 32'd5317, -32'd459, -32'd2418},
{-32'd1059, -32'd10330, 32'd7049, -32'd8816},
{-32'd4392, 32'd3643, 32'd2746, 32'd655},
{32'd4920, -32'd7565, -32'd6097, 32'd5892},
{-32'd2156, 32'd5244, -32'd2199, -32'd2112},
{-32'd3308, 32'd15383, -32'd10370, -32'd441},
{-32'd2574, 32'd4901, -32'd4147, 32'd5886},
{-32'd206, 32'd2919, -32'd4284, -32'd7201},
{32'd4662, 32'd5005, 32'd2992, 32'd1828},
{-32'd6460, 32'd2554, -32'd7194, -32'd6894},
{32'd4501, 32'd867, -32'd620, -32'd2071},
{-32'd7966, 32'd354, -32'd674, -32'd1047},
{-32'd10799, -32'd10875, -32'd1450, 32'd2928},
{-32'd10221, -32'd11392, 32'd13787, -32'd2936},
{32'd12701, 32'd9089, 32'd10842, -32'd2401},
{32'd5297, 32'd8388, 32'd2633, -32'd3888},
{-32'd14148, -32'd7211, -32'd2230, -32'd3695},
{-32'd8003, 32'd7844, 32'd5054, 32'd5099},
{32'd11547, -32'd4417, -32'd6354, 32'd1516},
{32'd3949, 32'd8141, 32'd10668, -32'd8112},
{32'd6365, -32'd898, 32'd3834, 32'd2421},
{32'd7816, -32'd266, -32'd1134, 32'd5689},
{32'd9415, 32'd11773, 32'd2219, 32'd3926},
{32'd1338, -32'd3753, 32'd3952, -32'd6833},
{-32'd6463, -32'd13767, 32'd2673, -32'd4013},
{-32'd3913, -32'd921, 32'd3244, -32'd273},
{32'd1758, 32'd4205, 32'd15470, -32'd4327},
{32'd10954, -32'd12347, 32'd5923, -32'd3597},
{32'd1534, -32'd10951, -32'd4396, -32'd5851},
{-32'd929, 32'd3887, -32'd6641, 32'd6706},
{-32'd7901, -32'd104, 32'd12145, 32'd1073},
{32'd2276, 32'd1894, 32'd3583, -32'd403},
{-32'd5976, -32'd2892, 32'd2287, 32'd2687},
{-32'd3481, 32'd14598, -32'd16347, -32'd2714},
{32'd254, 32'd6108, 32'd824, 32'd5244},
{-32'd5303, 32'd1151, -32'd2173, 32'd865},
{32'd3764, -32'd4231, -32'd7026, 32'd1838},
{-32'd4666, 32'd9645, -32'd7512, 32'd1871},
{-32'd7241, 32'd952, 32'd1441, -32'd2718},
{-32'd3544, -32'd4049, -32'd17283, 32'd7583},
{-32'd3223, 32'd10745, 32'd4804, -32'd7927},
{32'd325, -32'd1135, -32'd2528, 32'd2197},
{-32'd378, -32'd608, 32'd1251, -32'd5864},
{-32'd7835, 32'd4362, -32'd2374, 32'd4789},
{32'd756, 32'd4656, 32'd1723, 32'd4511},
{32'd3313, 32'd8251, -32'd7943, 32'd2764},
{32'd14217, 32'd10303, 32'd5458, 32'd5668},
{32'd1571, 32'd3303, -32'd3087, -32'd1130},
{-32'd2110, -32'd1485, -32'd7604, 32'd2021},
{-32'd4970, 32'd128, -32'd1184, 32'd1869},
{32'd8824, -32'd1581, -32'd11187, -32'd5616},
{32'd8721, -32'd2684, 32'd6732, -32'd2098},
{-32'd2301, -32'd5489, 32'd7610, 32'd13025},
{32'd6855, 32'd6165, 32'd2619, -32'd4239},
{32'd7133, 32'd5926, 32'd2628, 32'd12322},
{-32'd12977, -32'd8264, -32'd8609, -32'd9203},
{32'd5761, -32'd4920, -32'd3240, 32'd3840},
{-32'd8650, -32'd4268, -32'd14805, -32'd2664},
{-32'd6982, 32'd2862, -32'd6932, -32'd3564},
{-32'd818, 32'd11922, 32'd1694, 32'd835},
{-32'd3425, -32'd1919, -32'd257, 32'd585},
{32'd7078, 32'd11580, 32'd6759, 32'd1612},
{-32'd2658, 32'd1068, 32'd8754, -32'd208},
{-32'd12514, 32'd748, -32'd8817, 32'd8332},
{32'd138, -32'd8476, -32'd3163, -32'd349},
{-32'd15067, 32'd2185, -32'd5112, -32'd3212},
{32'd1830, -32'd245, 32'd5339, -32'd3025},
{32'd10122, 32'd3077, 32'd1630, -32'd1865},
{32'd6416, -32'd4288, -32'd17, -32'd2545},
{-32'd307, 32'd1696, -32'd4966, 32'd7271}
},
{{32'd412, -32'd1066, 32'd13054, -32'd12508},
{32'd8521, -32'd10301, -32'd1454, -32'd8063},
{-32'd8084, 32'd6262, 32'd6668, 32'd454},
{-32'd38, 32'd6901, 32'd7189, 32'd1013},
{-32'd1296, 32'd314, 32'd9377, 32'd91},
{-32'd2930, 32'd5124, -32'd6801, -32'd1235},
{32'd7162, -32'd412, 32'd4909, 32'd1700},
{32'd8400, 32'd1267, -32'd10308, -32'd7370},
{32'd10994, 32'd9198, 32'd5087, 32'd8587},
{32'd9501, 32'd8843, 32'd5727, 32'd175},
{-32'd6263, 32'd1638, -32'd140, 32'd10996},
{32'd3617, -32'd4716, -32'd3891, -32'd4768},
{-32'd13204, -32'd5145, 32'd5873, 32'd314},
{-32'd2440, -32'd4258, -32'd5422, 32'd3693},
{-32'd1026, -32'd988, -32'd5647, -32'd10989},
{-32'd4870, 32'd2633, -32'd2186, -32'd3060},
{32'd7346, 32'd2051, 32'd6380, -32'd13891},
{32'd7703, -32'd8706, 32'd1899, 32'd13890},
{-32'd10637, -32'd4299, -32'd6159, 32'd3860},
{-32'd9301, -32'd542, 32'd5084, -32'd2145},
{-32'd7549, -32'd1818, 32'd8993, 32'd3490},
{-32'd5627, -32'd5775, -32'd8139, 32'd552},
{-32'd1512, -32'd12715, 32'd5571, -32'd4877},
{-32'd5294, 32'd2391, 32'd5179, 32'd2396},
{32'd6856, 32'd6658, 32'd12251, -32'd432},
{-32'd2671, -32'd3541, 32'd2296, 32'd5818},
{32'd6366, -32'd14324, 32'd2245, -32'd1219},
{-32'd3018, -32'd8603, 32'd3463, 32'd7310},
{-32'd10612, 32'd11642, 32'd3393, 32'd6044},
{32'd771, 32'd3200, -32'd8382, 32'd3913},
{-32'd9078, -32'd11858, -32'd1212, -32'd1818},
{-32'd8066, -32'd12234, -32'd5674, -32'd3287},
{32'd8504, 32'd5443, 32'd6274, -32'd4452},
{-32'd6416, -32'd8614, -32'd1671, -32'd4574},
{32'd17030, 32'd5894, 32'd10060, 32'd3850},
{-32'd1398, 32'd10437, 32'd7173, 32'd14983},
{32'd2982, 32'd3962, -32'd8752, -32'd3859},
{32'd10141, 32'd1515, -32'd1318, -32'd6220},
{-32'd1324, -32'd3773, -32'd6671, -32'd7327},
{32'd15844, 32'd5207, 32'd2784, 32'd6616},
{-32'd6979, 32'd6464, -32'd6667, -32'd11212},
{32'd7386, -32'd2518, 32'd5036, 32'd6311},
{32'd6433, -32'd4531, -32'd1575, 32'd1811},
{-32'd8061, -32'd5838, -32'd2314, -32'd14839},
{-32'd1294, -32'd4204, 32'd1012, -32'd6169},
{32'd5814, -32'd3981, -32'd3569, 32'd10318},
{-32'd9656, -32'd4641, -32'd2918, 32'd1693},
{32'd5168, -32'd10485, -32'd6392, -32'd1799},
{-32'd706, 32'd4463, 32'd15495, 32'd1687},
{32'd3720, -32'd2747, 32'd6484, -32'd2048},
{-32'd3983, -32'd3551, 32'd7254, -32'd7909},
{32'd2435, 32'd485, 32'd4709, -32'd1414},
{-32'd4509, 32'd1970, -32'd1825, 32'd10615},
{-32'd3390, -32'd2612, 32'd8372, -32'd7858},
{32'd2515, 32'd4748, 32'd1357, -32'd13460},
{-32'd4609, -32'd1410, -32'd12793, -32'd2205},
{32'd9248, 32'd3828, 32'd13596, 32'd3334},
{-32'd6557, -32'd2604, -32'd7918, -32'd9626},
{-32'd14394, -32'd609, -32'd12617, -32'd9533},
{-32'd6446, -32'd6759, 32'd362, -32'd2027},
{32'd5829, -32'd9262, 32'd3606, 32'd11347},
{-32'd3041, 32'd656, 32'd505, -32'd339},
{-32'd5000, -32'd4175, -32'd4220, 32'd2282},
{-32'd8217, 32'd560, 32'd623, 32'd4033},
{32'd4048, 32'd5185, 32'd4050, -32'd1036},
{32'd9686, 32'd9705, 32'd13993, 32'd1392},
{32'd1979, -32'd5210, -32'd2981, 32'd6587},
{32'd3072, -32'd1771, -32'd1141, -32'd3066},
{-32'd3645, 32'd1814, 32'd2850, -32'd6432},
{32'd3185, 32'd7422, 32'd2295, 32'd6462},
{-32'd4172, 32'd3978, 32'd6401, -32'd6473},
{-32'd10267, 32'd7183, -32'd3338, -32'd5616},
{-32'd6191, 32'd4922, -32'd9663, -32'd9055},
{-32'd13405, -32'd1904, 32'd9115, 32'd4985},
{32'd1507, 32'd4528, 32'd5459, -32'd2960},
{32'd7383, 32'd11576, 32'd7380, -32'd14347},
{-32'd3580, -32'd7249, -32'd8808, -32'd1986},
{-32'd5115, -32'd10955, -32'd10486, 32'd9428},
{-32'd1591, 32'd10043, 32'd5636, 32'd1180},
{32'd14617, 32'd4522, 32'd1531, 32'd6229},
{32'd3082, -32'd4081, 32'd2035, -32'd4125},
{-32'd1434, 32'd4686, -32'd5714, 32'd446},
{-32'd6492, -32'd4838, -32'd4963, 32'd1379},
{32'd6944, -32'd6551, -32'd17533, -32'd4157},
{32'd4499, -32'd1601, -32'd9327, -32'd3086},
{-32'd12355, 32'd393, 32'd1109, 32'd7507},
{32'd1161, 32'd5980, 32'd9561, 32'd1359},
{-32'd11271, -32'd5788, 32'd1637, -32'd1401},
{-32'd64, -32'd9299, -32'd5959, -32'd8222},
{-32'd6557, -32'd4926, -32'd7188, -32'd4614},
{32'd8385, 32'd275, -32'd1007, 32'd3698},
{-32'd63, -32'd6162, 32'd440, -32'd2102},
{32'd14157, 32'd1147, 32'd6261, 32'd3012},
{32'd3805, -32'd5305, 32'd6175, -32'd2307},
{-32'd6084, 32'd3932, -32'd2018, -32'd3130},
{32'd1977, -32'd4428, -32'd13910, -32'd7775},
{32'd9694, 32'd10101, -32'd4506, -32'd3980},
{32'd5341, 32'd8081, 32'd2671, 32'd5813},
{32'd7166, 32'd1968, 32'd9291, 32'd2419},
{32'd8078, 32'd5982, -32'd3966, -32'd3250},
{-32'd3971, -32'd4325, -32'd11600, -32'd10001},
{-32'd2898, 32'd6186, 32'd6172, -32'd2351},
{-32'd950, 32'd281, -32'd14135, 32'd1223},
{32'd2276, 32'd5733, 32'd3988, -32'd5949},
{-32'd1883, 32'd11656, -32'd5216, 32'd5534},
{32'd8543, -32'd3753, 32'd817, 32'd5148},
{-32'd6135, -32'd8285, -32'd2859, 32'd7662},
{-32'd11904, 32'd3005, 32'd3930, -32'd9543},
{32'd17013, 32'd5900, -32'd3540, -32'd5064},
{32'd8608, 32'd3831, 32'd2172, 32'd3972},
{-32'd10622, 32'd4267, -32'd2864, -32'd7695},
{-32'd1557, 32'd3967, -32'd4503, -32'd5978},
{32'd807, -32'd2482, 32'd6745, 32'd3617},
{-32'd936, -32'd3298, 32'd10441, -32'd7079},
{-32'd1483, 32'd4181, -32'd1626, -32'd14768},
{32'd3348, -32'd2886, 32'd11460, 32'd5405},
{-32'd1012, 32'd2468, -32'd2920, -32'd5322},
{-32'd3512, 32'd1237, 32'd3007, 32'd2130},
{32'd10093, 32'd5390, 32'd11557, 32'd6973},
{32'd5544, 32'd11537, 32'd12034, 32'd8090},
{-32'd5858, 32'd8341, 32'd9530, -32'd5589},
{32'd9138, 32'd6962, 32'd12585, -32'd1446},
{32'd1745, -32'd14483, 32'd4590, 32'd7659},
{32'd3276, 32'd368, -32'd2967, 32'd4473},
{-32'd10136, -32'd5420, -32'd6077, 32'd3590},
{-32'd7245, 32'd4511, 32'd7012, -32'd5769},
{-32'd845, -32'd834, -32'd6235, 32'd9059},
{32'd281, 32'd5655, -32'd286, 32'd3281},
{32'd4420, -32'd5383, -32'd13666, -32'd10965},
{-32'd9766, 32'd1947, 32'd6467, -32'd1025},
{-32'd7770, 32'd2866, 32'd3534, 32'd12267},
{32'd9411, 32'd3648, -32'd5723, -32'd8262},
{-32'd121, -32'd11796, -32'd8777, 32'd2626},
{32'd2694, 32'd11080, 32'd1361, -32'd2666},
{32'd12090, -32'd676, 32'd4043, -32'd10590},
{32'd11051, 32'd3679, -32'd128, -32'd4599},
{-32'd3544, -32'd7706, 32'd1244, -32'd5755},
{32'd3259, -32'd8545, -32'd2208, -32'd3082},
{32'd2510, -32'd1871, 32'd3601, 32'd4334},
{-32'd941, -32'd10466, -32'd14970, -32'd7109},
{-32'd3888, -32'd2137, 32'd1535, 32'd1058},
{-32'd10206, -32'd2383, -32'd19039, 32'd2842},
{-32'd2637, 32'd1393, 32'd7473, 32'd2210},
{-32'd9382, -32'd835, -32'd904, -32'd1672},
{32'd7793, -32'd1483, 32'd8881, -32'd4841},
{32'd2596, -32'd2688, 32'd933, 32'd745},
{32'd13920, -32'd3190, -32'd1181, -32'd2120},
{-32'd8169, 32'd4706, 32'd2450, 32'd4504},
{32'd4499, 32'd3727, 32'd9318, -32'd699},
{-32'd2144, -32'd9808, -32'd9777, 32'd390},
{-32'd7636, -32'd8931, -32'd9391, -32'd3659},
{32'd15057, 32'd5751, 32'd504, 32'd7946},
{-32'd8439, 32'd940, -32'd3121, 32'd3602},
{-32'd5434, 32'd1715, -32'd10399, -32'd5864},
{-32'd8985, -32'd6188, -32'd12124, 32'd2222},
{32'd15973, -32'd1149, 32'd6585, -32'd951},
{32'd5584, -32'd3550, -32'd3591, 32'd9787},
{-32'd8619, -32'd5602, 32'd3170, -32'd2303},
{32'd2068, -32'd8735, 32'd2993, 32'd7429},
{-32'd4093, 32'd2642, -32'd4863, -32'd1929},
{-32'd922, 32'd61, 32'd156, -32'd6795},
{32'd2949, 32'd6482, 32'd2574, -32'd13564},
{-32'd1661, -32'd1180, 32'd2823, -32'd7843},
{32'd813, -32'd4116, 32'd11346, -32'd3856},
{-32'd4494, 32'd13969, -32'd554, 32'd7497},
{-32'd8890, -32'd4770, 32'd1842, -32'd3750},
{32'd12844, -32'd537, -32'd2264, -32'd1974},
{-32'd3397, -32'd1986, 32'd2356, -32'd9315},
{32'd1306, -32'd2589, -32'd8962, -32'd4267},
{-32'd6134, 32'd1204, -32'd7279, -32'd2122},
{-32'd4521, -32'd1740, -32'd11300, 32'd9014},
{-32'd285, 32'd4806, -32'd11694, 32'd8483},
{32'd11269, 32'd4163, 32'd8567, 32'd9854},
{-32'd9831, 32'd125, 32'd4679, 32'd8076},
{-32'd1515, 32'd1685, 32'd4489, 32'd2549},
{32'd1072, 32'd2521, -32'd3855, -32'd9892},
{32'd13842, 32'd9786, -32'd898, -32'd739},
{-32'd3766, 32'd3942, 32'd3796, 32'd5329},
{32'd13995, 32'd6867, 32'd8408, 32'd3689},
{-32'd5194, -32'd9105, -32'd2406, -32'd11970},
{-32'd3120, -32'd3139, -32'd5041, 32'd6458},
{-32'd3167, -32'd4439, -32'd1315, -32'd6228},
{-32'd3592, -32'd11781, -32'd3855, 32'd9549},
{32'd2713, 32'd13119, -32'd76, -32'd7447},
{-32'd5967, 32'd3300, -32'd4944, 32'd872},
{-32'd232, -32'd541, -32'd253, -32'd7947},
{-32'd1559, 32'd4317, 32'd6875, 32'd5443},
{32'd16990, 32'd9606, -32'd329, 32'd3598},
{-32'd216, -32'd8240, 32'd364, 32'd1377},
{-32'd9764, 32'd4572, -32'd784, -32'd497},
{32'd9639, 32'd2661, 32'd7098, 32'd15810},
{-32'd6303, -32'd2702, -32'd3000, 32'd2360},
{32'd4320, 32'd794, -32'd15211, 32'd3457},
{32'd1421, -32'd4400, 32'd11206, 32'd9058},
{32'd6742, 32'd4207, -32'd1975, -32'd3495},
{32'd3277, -32'd2766, 32'd4780, -32'd4696},
{32'd9413, -32'd2825, 32'd3892, -32'd3436},
{-32'd1221, 32'd7909, 32'd13041, -32'd860},
{-32'd252, -32'd3706, 32'd4662, 32'd2783},
{32'd5694, -32'd3725, 32'd7, -32'd9586},
{-32'd12655, -32'd3376, -32'd7003, -32'd5510},
{-32'd1536, 32'd6839, 32'd2461, 32'd799},
{-32'd10583, -32'd7311, 32'd5850, 32'd4429},
{32'd9296, -32'd4871, 32'd2191, -32'd467},
{-32'd5828, -32'd6170, -32'd21270, -32'd1045},
{32'd865, 32'd1249, -32'd9806, 32'd4018},
{32'd5818, 32'd230, -32'd9031, 32'd3710},
{-32'd9997, -32'd2893, -32'd11945, -32'd990},
{-32'd3832, -32'd266, -32'd2386, 32'd5843},
{32'd7199, 32'd7325, -32'd1668, -32'd10664},
{32'd1523, 32'd1351, -32'd390, 32'd1408},
{32'd5676, -32'd3865, -32'd3536, -32'd6044},
{-32'd4818, -32'd2933, -32'd2254, 32'd1828},
{32'd7894, -32'd2414, 32'd1777, -32'd918},
{-32'd2936, -32'd4550, 32'd4906, -32'd1596},
{-32'd10302, -32'd14264, 32'd3462, -32'd8193},
{32'd2861, 32'd2951, 32'd14409, 32'd7417},
{-32'd8583, -32'd3184, -32'd5250, -32'd3550},
{32'd12376, 32'd2624, 32'd6482, -32'd5444},
{32'd753, -32'd9498, 32'd2618, -32'd6141},
{-32'd5341, -32'd10328, -32'd1931, 32'd2236},
{32'd4875, 32'd12095, 32'd5784, 32'd5631},
{32'd2866, 32'd5902, 32'd6988, 32'd1374},
{-32'd5615, 32'd2632, 32'd4333, -32'd2712},
{32'd938, -32'd3454, -32'd2504, 32'd722},
{32'd7560, 32'd919, 32'd7351, -32'd2105},
{32'd3501, -32'd4309, -32'd13351, 32'd2746},
{-32'd2631, -32'd3787, 32'd2396, -32'd6020},
{32'd4038, -32'd2739, 32'd7083, 32'd6449},
{-32'd984, 32'd3536, 32'd9290, -32'd4435},
{-32'd2418, -32'd12434, -32'd4029, 32'd5832},
{32'd563, 32'd5930, 32'd144, 32'd194},
{-32'd8680, 32'd3647, 32'd5651, 32'd15050},
{-32'd907, -32'd2717, 32'd969, -32'd9092},
{-32'd3359, -32'd7229, -32'd9523, -32'd1075},
{-32'd5486, 32'd3380, -32'd8040, -32'd1451},
{-32'd2545, 32'd3021, 32'd1567, -32'd9421},
{-32'd3859, 32'd3045, 32'd7672, 32'd11163},
{32'd5765, 32'd6007, -32'd1700, 32'd1368},
{-32'd12020, -32'd3408, -32'd3131, 32'd1639},
{-32'd8082, 32'd2494, 32'd9288, 32'd6844},
{-32'd3302, -32'd830, -32'd3774, 32'd2119},
{-32'd5847, -32'd4205, -32'd10799, -32'd3687},
{-32'd2571, 32'd7891, 32'd6261, 32'd11985},
{32'd3308, 32'd8703, -32'd206, -32'd326},
{32'd4417, -32'd3003, -32'd4706, -32'd2837},
{32'd4433, -32'd10773, -32'd7971, 32'd104},
{-32'd3118, 32'd2772, 32'd1049, 32'd469},
{32'd983, 32'd3653, -32'd7662, -32'd7786},
{32'd4212, 32'd6325, -32'd7790, -32'd5022},
{32'd1166, -32'd10584, -32'd3679, 32'd5101},
{-32'd7102, -32'd2990, -32'd3658, -32'd5444},
{32'd5438, 32'd4801, 32'd1967, -32'd3649},
{-32'd226, -32'd1263, 32'd919, -32'd568},
{-32'd5645, -32'd417, -32'd1700, -32'd3652},
{32'd8622, -32'd1326, 32'd14324, -32'd13},
{-32'd14420, 32'd1443, -32'd2239, 32'd5392},
{32'd8377, 32'd3024, 32'd1547, -32'd5772},
{-32'd5432, -32'd889, -32'd5651, -32'd472},
{-32'd2424, 32'd4024, 32'd9104, -32'd1953},
{-32'd2340, 32'd7612, 32'd7129, 32'd8791},
{32'd1914, -32'd4276, 32'd3813, -32'd10225},
{-32'd9585, -32'd8341, -32'd8265, 32'd6044},
{-32'd2918, 32'd1660, -32'd2111, 32'd316},
{-32'd6184, -32'd10898, 32'd4133, 32'd9392},
{32'd3950, 32'd7038, 32'd10167, 32'd818},
{-32'd5001, 32'd6611, -32'd971, -32'd651},
{-32'd3259, -32'd2158, 32'd3331, 32'd10085},
{-32'd10892, 32'd4533, -32'd6874, -32'd3896},
{-32'd3339, -32'd12111, 32'd2111, -32'd3236},
{-32'd6402, 32'd7193, 32'd6183, 32'd4261},
{32'd12354, -32'd4579, 32'd4927, -32'd7288},
{-32'd7273, 32'd875, 32'd2325, 32'd768},
{32'd6806, -32'd1680, -32'd9512, 32'd5689},
{32'd543, -32'd1793, -32'd2971, -32'd3056},
{-32'd4504, -32'd11560, 32'd4335, 32'd2065},
{32'd13216, 32'd8047, 32'd7759, 32'd2912},
{-32'd2301, 32'd1222, -32'd689, 32'd3660},
{32'd2973, -32'd7541, -32'd17735, -32'd8549},
{32'd2432, -32'd10792, -32'd8906, -32'd5197},
{32'd1184, 32'd3788, -32'd4158, -32'd18},
{32'd4772, 32'd7757, 32'd11108, 32'd487},
{-32'd1807, 32'd1313, -32'd1627, -32'd3607},
{-32'd2752, -32'd4447, 32'd9332, 32'd9225},
{32'd7486, 32'd8815, 32'd10046, -32'd3324},
{-32'd10536, -32'd10759, -32'd5403, 32'd524},
{32'd1334, 32'd8911, 32'd4532, 32'd1921},
{-32'd2569, 32'd1003, -32'd5610, -32'd1868},
{32'd12050, -32'd15841, 32'd1146, -32'd2299},
{32'd3285, -32'd322, -32'd2498, -32'd5985},
{-32'd9358, -32'd6088, 32'd14576, 32'd5893},
{32'd1956, 32'd7174, 32'd6249, 32'd3548},
{32'd3510, -32'd1254, -32'd1800, -32'd6},
{-32'd12376, 32'd3698, -32'd6824, -32'd7233},
{32'd10261, -32'd97, -32'd3906, 32'd821},
{32'd13021, -32'd2788, 32'd2513, -32'd11268},
{-32'd6742, -32'd72, -32'd108, 32'd3736},
{32'd1162, 32'd9868, -32'd4996, -32'd9249},
{32'd9879, -32'd1636, 32'd8244, 32'd4134},
{-32'd7681, 32'd1299, 32'd4110, 32'd7173}
},
{{32'd11841, 32'd3071, 32'd389, -32'd5691},
{-32'd16349, -32'd3457, 32'd2228, -32'd4448},
{32'd10128, 32'd8925, 32'd8211, 32'd9022},
{32'd15355, 32'd2373, 32'd12072, 32'd1020},
{-32'd7344, -32'd10828, -32'd4119, -32'd4574},
{-32'd2368, -32'd11497, -32'd2046, 32'd4586},
{32'd2551, 32'd8750, 32'd1380, 32'd9376},
{32'd1571, 32'd1650, 32'd9912, -32'd131},
{-32'd3219, 32'd8656, 32'd11678, 32'd10024},
{32'd8684, 32'd13213, 32'd8254, 32'd7023},
{-32'd3901, 32'd4500, -32'd5303, 32'd5843},
{32'd5386, -32'd4752, 32'd7193, 32'd9667},
{32'd2869, -32'd7194, 32'd6790, -32'd1888},
{32'd8563, -32'd10446, 32'd6035, 32'd1245},
{-32'd6967, -32'd10381, 32'd1698, 32'd1026},
{-32'd11911, -32'd11366, -32'd8745, -32'd4670},
{32'd14793, 32'd1957, 32'd4082, -32'd9562},
{-32'd8369, 32'd4746, 32'd14714, 32'd3665},
{32'd8047, -32'd9259, 32'd501, 32'd9725},
{-32'd8423, 32'd5911, -32'd8211, -32'd6233},
{32'd939, -32'd1732, -32'd3447, -32'd6091},
{-32'd12997, -32'd7280, -32'd2762, -32'd12602},
{-32'd16885, -32'd10245, 32'd4515, -32'd7204},
{32'd2120, -32'd11432, -32'd11218, -32'd10092},
{32'd3638, 32'd11324, 32'd2581, -32'd3591},
{32'd11895, 32'd1953, 32'd10430, -32'd2089},
{-32'd22743, 32'd5684, -32'd7398, -32'd7250},
{32'd1208, 32'd7375, 32'd12369, -32'd1110},
{32'd4914, -32'd6960, 32'd7862, -32'd1066},
{32'd8221, 32'd3262, 32'd1654, 32'd12420},
{-32'd11071, 32'd3155, -32'd712, -32'd6173},
{-32'd8178, -32'd10413, -32'd1222, -32'd7492},
{32'd5292, 32'd6401, 32'd6166, 32'd7047},
{32'd530, -32'd2941, 32'd4233, -32'd7414},
{32'd4055, 32'd15476, 32'd2175, 32'd8952},
{-32'd2433, 32'd7790, -32'd14341, -32'd1974},
{32'd8686, -32'd3142, 32'd9621, -32'd3751},
{32'd3595, -32'd11107, 32'd15262, -32'd20338},
{-32'd49, 32'd3217, 32'd2656, 32'd413},
{32'd12259, -32'd709, -32'd5029, 32'd3002},
{-32'd7544, 32'd1277, 32'd6435, -32'd14578},
{32'd4542, 32'd12651, -32'd3732, 32'd14756},
{-32'd4285, 32'd7079, -32'd7025, -32'd3802},
{32'd302, 32'd5549, -32'd2571, -32'd6871},
{-32'd6155, -32'd6502, -32'd3673, -32'd1286},
{32'd2900, 32'd11814, 32'd295, -32'd15125},
{-32'd3422, -32'd958, -32'd9866, -32'd11769},
{-32'd10642, -32'd6128, 32'd588, -32'd4996},
{-32'd10789, -32'd2415, 32'd6351, 32'd18273},
{-32'd21560, -32'd368, -32'd4957, 32'd2475},
{-32'd8314, -32'd4248, -32'd681, -32'd4086},
{32'd2049, -32'd2600, 32'd5779, 32'd1169},
{-32'd17831, 32'd449, -32'd10504, 32'd3925},
{32'd2418, -32'd9783, -32'd2644, -32'd7465},
{32'd834, 32'd6026, 32'd8181, 32'd614},
{-32'd3988, -32'd8143, -32'd3278, -32'd4884},
{32'd4414, 32'd5623, 32'd1670, 32'd5284},
{-32'd986, -32'd9999, 32'd3889, -32'd18},
{-32'd6492, -32'd4574, -32'd2444, -32'd2812},
{-32'd6171, -32'd5570, -32'd11222, 32'd6605},
{32'd9050, -32'd3644, 32'd4710, -32'd1911},
{32'd10844, 32'd2391, 32'd7248, -32'd1401},
{-32'd6713, -32'd6214, -32'd17279, -32'd3447},
{32'd3185, 32'd7838, -32'd447, 32'd1906},
{32'd4358, -32'd7399, -32'd784, 32'd6108},
{-32'd6656, 32'd7221, 32'd397, 32'd2365},
{32'd5638, 32'd1816, 32'd6031, -32'd9416},
{-32'd5233, -32'd212, -32'd5686, -32'd1456},
{-32'd6834, 32'd3984, 32'd9179, -32'd2023},
{32'd10941, 32'd5530, -32'd11733, -32'd484},
{-32'd18083, -32'd1203, -32'd9179, -32'd7159},
{-32'd2128, 32'd11957, 32'd8615, -32'd3023},
{-32'd2645, -32'd4137, 32'd5023, 32'd5437},
{32'd2589, 32'd2259, -32'd10032, -32'd761},
{-32'd276, -32'd858, 32'd6001, 32'd9321},
{32'd6552, 32'd6059, -32'd8076, -32'd7295},
{32'd11121, -32'd19474, -32'd3006, -32'd5232},
{32'd16360, -32'd5293, 32'd976, 32'd10957},
{32'd7699, 32'd9696, 32'd10954, -32'd3423},
{32'd10980, 32'd6234, -32'd5530, -32'd9108},
{-32'd2648, 32'd10561, 32'd12713, 32'd4966},
{32'd175, 32'd2809, -32'd4588, -32'd608},
{32'd367, 32'd316, -32'd6156, 32'd824},
{32'd8140, -32'd6624, -32'd4063, -32'd1719},
{32'd4713, 32'd1529, -32'd7554, -32'd1798},
{-32'd2646, -32'd2956, 32'd4917, -32'd3032},
{-32'd3234, 32'd3015, 32'd958, 32'd138},
{-32'd153, -32'd2444, -32'd9721, -32'd8701},
{-32'd6450, -32'd13935, 32'd10521, -32'd2355},
{-32'd18983, -32'd1131, 32'd2559, 32'd8402},
{32'd5844, 32'd7862, 32'd13668, 32'd5249},
{-32'd19203, 32'd1781, 32'd289, 32'd1429},
{-32'd5700, 32'd5915, 32'd2758, 32'd5},
{32'd9120, 32'd5323, 32'd3448, -32'd5475},
{-32'd6363, 32'd5547, 32'd11941, 32'd11303},
{32'd1585, -32'd2287, 32'd4290, -32'd8805},
{32'd5772, 32'd10995, 32'd870, 32'd6886},
{-32'd2714, 32'd5759, -32'd330, 32'd12585},
{32'd12937, -32'd3960, 32'd5244, 32'd13348},
{-32'd4498, 32'd468, 32'd6001, 32'd881},
{-32'd12792, -32'd13367, -32'd12194, -32'd19078},
{-32'd15103, 32'd4916, -32'd7244, -32'd6788},
{32'd26292, -32'd10514, -32'd3983, -32'd5592},
{32'd2320, 32'd4060, -32'd5932, 32'd994},
{-32'd6013, 32'd4628, -32'd2952, -32'd9248},
{-32'd884, 32'd979, -32'd8042, -32'd4001},
{-32'd3669, -32'd5029, 32'd8793, 32'd1069},
{32'd2281, 32'd8539, 32'd6452, -32'd7771},
{32'd5548, 32'd5773, -32'd5292, -32'd648},
{-32'd3138, -32'd533, -32'd13280, -32'd9697},
{-32'd1899, 32'd2147, -32'd12774, -32'd10343},
{32'd17326, -32'd11545, -32'd13746, -32'd1835},
{32'd11709, 32'd11958, 32'd14130, 32'd8835},
{-32'd1997, 32'd7928, 32'd3676, -32'd4977},
{-32'd7096, -32'd6826, -32'd4423, -32'd5038},
{-32'd22392, -32'd2626, -32'd1793, -32'd4759},
{-32'd9937, 32'd13280, -32'd7347, -32'd1007},
{-32'd3226, 32'd8275, -32'd4078, 32'd1018},
{32'd474, 32'd3385, -32'd4248, 32'd2928},
{-32'd11528, 32'd17825, 32'd5058, 32'd5257},
{32'd1815, -32'd6024, 32'd5258, 32'd3282},
{32'd5072, -32'd9515, 32'd1584, -32'd601},
{-32'd1342, -32'd992, 32'd8804, -32'd1093},
{-32'd6304, -32'd10877, 32'd3065, 32'd237},
{32'd2699, -32'd19140, 32'd1042, 32'd12495},
{32'd8700, 32'd166, 32'd3364, 32'd16609},
{32'd6396, -32'd8499, -32'd9831, 32'd4674},
{32'd2600, 32'd1707, -32'd3015, -32'd604},
{-32'd1938, -32'd9886, -32'd7847, -32'd5935},
{32'd8642, -32'd2578, -32'd5965, -32'd3630},
{-32'd13765, 32'd7314, -32'd6698, 32'd1880},
{32'd1762, -32'd2496, -32'd10061, -32'd2700},
{-32'd908, -32'd10976, -32'd7838, -32'd9839},
{-32'd8361, -32'd2384, -32'd4510, 32'd562},
{32'd4477, 32'd4416, 32'd10229, -32'd3544},
{-32'd7980, 32'd5236, 32'd2227, 32'd1250},
{-32'd2525, 32'd15, 32'd4239, -32'd14002},
{32'd9433, 32'd1359, -32'd269, -32'd2436},
{32'd4910, -32'd6889, 32'd15786, 32'd8744},
{-32'd8690, 32'd13, -32'd14205, -32'd14241},
{-32'd1589, 32'd4212, -32'd22368, -32'd8850},
{32'd333, -32'd5872, -32'd9534, -32'd7684},
{-32'd6564, -32'd8664, 32'd8731, 32'd4817},
{-32'd16542, -32'd3169, 32'd12579, -32'd314},
{32'd8223, 32'd7518, -32'd9926, -32'd2098},
{-32'd3221, 32'd10071, 32'd12063, 32'd6171},
{-32'd11363, -32'd3836, 32'd2199, 32'd1022},
{-32'd864, -32'd531, -32'd7226, -32'd5503},
{-32'd3803, 32'd1247, 32'd6717, 32'd8901},
{32'd2361, -32'd11952, -32'd3211, 32'd1777},
{32'd8017, -32'd7425, -32'd1522, -32'd8551},
{32'd11629, -32'd2050, 32'd6552, 32'd12203},
{-32'd10605, -32'd5612, -32'd2137, -32'd9266},
{-32'd712, 32'd7924, 32'd4, -32'd13609},
{-32'd5471, 32'd7057, 32'd3710, -32'd1459},
{32'd783, -32'd7314, 32'd8090, -32'd4579},
{32'd11481, 32'd13218, 32'd7581, 32'd12104},
{32'd5918, 32'd9206, 32'd9743, 32'd10684},
{-32'd10030, -32'd10682, -32'd4738, -32'd8438},
{32'd3175, 32'd757, 32'd2687, 32'd7365},
{-32'd2202, 32'd3975, -32'd10528, 32'd5647},
{-32'd335, -32'd716, -32'd1314, 32'd568},
{-32'd10317, -32'd3565, -32'd11439, -32'd7318},
{32'd9763, -32'd8138, 32'd2293, 32'd582},
{-32'd6572, -32'd3896, -32'd4406, 32'd4766},
{32'd6051, 32'd2286, -32'd3542, 32'd8137},
{-32'd7504, 32'd2949, -32'd8103, 32'd2451},
{32'd2459, -32'd3249, -32'd10268, -32'd5232},
{32'd11089, -32'd21535, -32'd4652, -32'd16767},
{32'd218, -32'd6802, -32'd7306, -32'd3529},
{-32'd869, -32'd1738, 32'd64, 32'd10249},
{32'd9128, 32'd4713, -32'd7894, 32'd5637},
{32'd11321, 32'd10876, 32'd11277, 32'd11821},
{32'd8574, -32'd7283, -32'd1169, -32'd7600},
{32'd3789, -32'd6509, 32'd13282, 32'd4846},
{-32'd289, -32'd4480, -32'd6803, -32'd443},
{32'd10058, -32'd4935, 32'd1151, 32'd8225},
{-32'd7234, -32'd9761, 32'd8054, -32'd5530},
{32'd4324, -32'd4379, -32'd14254, 32'd1528},
{-32'd12643, -32'd6381, 32'd3607, -32'd6607},
{-32'd4173, -32'd4809, -32'd6733, -32'd15087},
{-32'd6302, -32'd6397, -32'd9592, -32'd4925},
{32'd5288, -32'd10999, -32'd10269, -32'd2598},
{32'd2894, -32'd9849, -32'd10138, 32'd936},
{-32'd2898, -32'd87, -32'd6208, -32'd9207},
{-32'd55, -32'd216, 32'd11234, 32'd4678},
{-32'd5262, 32'd6536, 32'd9138, 32'd12307},
{-32'd5598, 32'd2873, -32'd2622, 32'd4164},
{32'd8385, -32'd3160, 32'd5985, 32'd2194},
{-32'd3988, -32'd6427, 32'd2016, 32'd2761},
{-32'd5326, -32'd5049, 32'd5560, -32'd3114},
{32'd4517, -32'd8744, -32'd85, -32'd8774},
{-32'd1039, -32'd3221, 32'd6705, 32'd10150},
{32'd1552, -32'd5781, 32'd3757, 32'd7784},
{-32'd1080, 32'd10720, -32'd4376, 32'd3037},
{-32'd6314, 32'd301, -32'd388, -32'd346},
{32'd957, 32'd2951, -32'd2410, -32'd11862},
{-32'd7821, 32'd3653, -32'd5452, -32'd9139},
{32'd1170, -32'd236, 32'd7425, 32'd16091},
{-32'd10345, 32'd3232, -32'd225, -32'd3602},
{-32'd11111, -32'd14615, -32'd7634, -32'd8016},
{-32'd7258, 32'd6638, 32'd1728, -32'd11942},
{32'd929, 32'd3531, -32'd3987, -32'd2797},
{32'd21536, -32'd2802, 32'd5506, 32'd8946},
{32'd3292, -32'd10184, -32'd6783, -32'd7010},
{32'd15962, -32'd2514, -32'd694, 32'd320},
{32'd3200, -32'd955, -32'd98, 32'd7549},
{-32'd1967, -32'd14008, -32'd5119, -32'd8614},
{32'd768, 32'd2214, 32'd20076, 32'd8594},
{32'd5661, -32'd1358, 32'd8419, 32'd2659},
{-32'd10150, 32'd1943, -32'd272, -32'd3069},
{-32'd15274, 32'd5520, -32'd1042, -32'd10442},
{-32'd683, -32'd9413, -32'd1557, 32'd12508},
{32'd15312, -32'd5213, 32'd22126, 32'd609},
{-32'd5448, -32'd813, -32'd4917, -32'd10615},
{-32'd2619, -32'd2770, -32'd1030, -32'd6258},
{32'd8319, 32'd11443, -32'd2844, 32'd6260},
{-32'd7825, 32'd2394, 32'd7786, -32'd2839},
{32'd17088, 32'd12885, 32'd2380, 32'd3664},
{-32'd2248, 32'd8029, 32'd2637, 32'd3572},
{-32'd2895, -32'd4088, -32'd5598, 32'd2038},
{-32'd3037, 32'd8824, -32'd9182, -32'd3453},
{32'd905, 32'd4500, 32'd10313, 32'd12069},
{-32'd5634, -32'd3376, 32'd10022, -32'd1320},
{-32'd295, -32'd12917, -32'd13510, 32'd7139},
{32'd11196, -32'd506, -32'd8850, -32'd816},
{32'd12124, -32'd51, 32'd2532, 32'd2614},
{-32'd5634, 32'd219, -32'd10642, -32'd4835},
{32'd15784, -32'd2573, -32'd3418, -32'd795},
{32'd4434, 32'd7399, 32'd1905, -32'd1385},
{-32'd8261, -32'd4837, -32'd1421, -32'd12880},
{-32'd13473, 32'd32, 32'd3441, -32'd3676},
{-32'd1049, 32'd7088, 32'd3180, 32'd5913},
{-32'd12100, -32'd8, -32'd7806, -32'd4021},
{32'd1446, -32'd9839, 32'd1662, -32'd3826},
{-32'd1672, -32'd556, -32'd4908, -32'd6391},
{-32'd20565, -32'd6576, 32'd4003, -32'd3362},
{-32'd6978, 32'd4565, 32'd15540, -32'd9763},
{32'd7143, 32'd8522, 32'd249, 32'd5604},
{-32'd3700, 32'd9115, 32'd7367, 32'd9573},
{-32'd7795, 32'd6308, -32'd10409, -32'd2466},
{-32'd1985, -32'd7453, 32'd6488, 32'd1161},
{-32'd5434, -32'd2934, -32'd6116, -32'd10983},
{-32'd9536, 32'd2265, -32'd4790, -32'd2420},
{32'd8581, 32'd8803, 32'd9796, 32'd9631},
{32'd17985, -32'd6254, -32'd8074, -32'd2745},
{32'd2719, -32'd1868, 32'd5131, 32'd1963},
{-32'd10157, 32'd15590, -32'd1622, 32'd8005},
{32'd1348, -32'd7385, 32'd6673, 32'd12745},
{32'd4698, -32'd1556, 32'd2753, -32'd18356},
{-32'd10279, 32'd457, -32'd13555, 32'd508},
{-32'd5475, 32'd4410, 32'd8491, 32'd15588},
{-32'd7568, -32'd1880, 32'd7379, 32'd2300},
{32'd4631, 32'd1219, -32'd11393, -32'd12976},
{-32'd1375, -32'd2177, -32'd5756, -32'd902},
{32'd3978, -32'd3497, -32'd688, -32'd3307},
{-32'd1549, -32'd7594, -32'd7576, -32'd4706},
{32'd7132, -32'd4149, -32'd11190, -32'd3663},
{-32'd5502, -32'd13477, -32'd13750, -32'd7125},
{32'd498, 32'd2253, 32'd413, -32'd2855},
{-32'd7060, 32'd8160, 32'd13859, 32'd10504},
{32'd154, -32'd624, -32'd3894, -32'd9734},
{-32'd1944, -32'd5638, 32'd411, -32'd1866},
{-32'd2914, -32'd6101, -32'd3590, -32'd1014},
{-32'd16523, -32'd594, 32'd3399, -32'd2063},
{-32'd21341, 32'd6710, 32'd1294, 32'd3536},
{32'd14327, 32'd9659, 32'd4615, 32'd10907},
{-32'd7877, 32'd4883, 32'd408, 32'd10925},
{-32'd12080, -32'd1536, -32'd2622, 32'd6651},
{-32'd13563, -32'd3732, 32'd2267, 32'd5876},
{32'd5858, 32'd10941, -32'd1214, -32'd9939},
{32'd660, 32'd11665, 32'd9600, 32'd20186},
{-32'd8397, -32'd2733, -32'd3777, -32'd427},
{-32'd11165, 32'd8940, -32'd2712, -32'd3599},
{-32'd2923, -32'd2112, -32'd4057, -32'd1669},
{32'd5783, -32'd1323, -32'd2348, -32'd8568},
{32'd11048, 32'd12539, 32'd8469, 32'd11148},
{-32'd4808, 32'd54, 32'd9348, -32'd1981},
{-32'd4869, -32'd11218, -32'd152, -32'd897},
{32'd2970, -32'd6574, 32'd4256, -32'd3450},
{32'd298, 32'd5874, 32'd7431, 32'd8964},
{-32'd1716, 32'd8634, 32'd2060, 32'd4217},
{32'd9735, 32'd6619, -32'd705, -32'd2151},
{32'd10082, -32'd5997, -32'd13381, 32'd5056},
{32'd5070, 32'd17357, 32'd18058, 32'd13838},
{-32'd7389, -32'd6588, -32'd2316, -32'd4422},
{-32'd9312, 32'd4844, -32'd11740, -32'd1061},
{-32'd468, -32'd3533, -32'd6005, 32'd1105},
{32'd11264, -32'd4686, 32'd4916, -32'd1942},
{32'd13544, -32'd5610, -32'd900, -32'd1431},
{32'd4731, 32'd3589, -32'd4319, 32'd6058},
{32'd7300, 32'd4810, 32'd2141, 32'd15079},
{-32'd22, -32'd10656, -32'd8157, -32'd8855},
{-32'd13501, -32'd885, -32'd4334, 32'd5780},
{-32'd10546, 32'd2161, 32'd1661, -32'd9136},
{32'd6739, -32'd6111, 32'd4247, -32'd5325},
{32'd4482, 32'd1154, 32'd2896, 32'd5124},
{-32'd459, 32'd6546, 32'd4263, 32'd5540},
{-32'd922, 32'd8866, -32'd7651, 32'd9259},
{-32'd15828, -32'd5909, -32'd2818, -32'd6726}
},
{{-32'd4192, -32'd650, -32'd4095, 32'd8525},
{32'd15007, -32'd787, -32'd5527, -32'd11863},
{32'd8135, 32'd9337, 32'd2091, -32'd16218},
{-32'd8048, -32'd11434, -32'd500, -32'd527},
{32'd3402, 32'd12111, 32'd6913, -32'd8755},
{32'd16, 32'd3519, -32'd3194, -32'd3685},
{-32'd2167, 32'd6632, -32'd165, -32'd3312},
{32'd2318, 32'd3657, -32'd9033, -32'd2197},
{-32'd5342, 32'd11657, -32'd6412, 32'd7646},
{32'd9519, -32'd583, 32'd3127, 32'd233},
{-32'd11037, -32'd927, -32'd3351, 32'd6932},
{-32'd5044, 32'd1793, -32'd990, 32'd4369},
{-32'd1042, -32'd531, -32'd2257, -32'd3491},
{-32'd6411, -32'd9560, 32'd3965, 32'd3019},
{-32'd15334, -32'd2801, -32'd8880, -32'd502},
{-32'd9982, -32'd3348, 32'd11160, 32'd5536},
{32'd1964, -32'd3379, -32'd1627, 32'd843},
{32'd7689, 32'd5394, 32'd3013, 32'd85},
{-32'd5753, 32'd3881, -32'd2139, -32'd1944},
{-32'd7652, 32'd1077, 32'd7143, 32'd5872},
{32'd1277, 32'd2207, -32'd166, -32'd4885},
{32'd1545, 32'd5472, -32'd3827, 32'd12899},
{32'd7427, -32'd4275, -32'd4623, 32'd6441},
{-32'd10950, -32'd7136, -32'd3540, 32'd433},
{32'd3204, -32'd9958, 32'd14734, -32'd6165},
{32'd5553, -32'd9392, -32'd7770, -32'd4569},
{-32'd2833, -32'd172, -32'd4465, 32'd10649},
{32'd5124, 32'd332, 32'd13706, 32'd6838},
{32'd8235, 32'd12175, 32'd8728, -32'd5967},
{-32'd12233, 32'd9328, 32'd4851, -32'd4228},
{-32'd5704, -32'd154, -32'd6132, -32'd3149},
{-32'd611, 32'd2115, -32'd4024, 32'd5232},
{-32'd540, 32'd3078, -32'd3219, 32'd8938},
{32'd649, -32'd9263, 32'd5957, -32'd300},
{32'd15372, 32'd6830, 32'd8848, 32'd5786},
{32'd202, 32'd2601, -32'd13068, 32'd203},
{32'd7227, 32'd13558, 32'd11396, -32'd2571},
{32'd6821, -32'd6935, 32'd4523, -32'd11432},
{-32'd13347, -32'd5695, -32'd2721, 32'd5497},
{-32'd4138, 32'd7363, 32'd3867, 32'd8496},
{32'd13390, -32'd8407, 32'd11355, -32'd11855},
{-32'd6577, 32'd16139, -32'd2780, 32'd5163},
{-32'd13547, -32'd1099, 32'd18890, 32'd11903},
{-32'd5267, -32'd22278, 32'd2435, -32'd1674},
{-32'd15395, -32'd432, -32'd2935, 32'd1962},
{-32'd7338, -32'd14137, 32'd2528, -32'd654},
{-32'd8449, -32'd413, -32'd8634, -32'd9038},
{-32'd14413, -32'd7825, 32'd3549, -32'd11825},
{-32'd7653, 32'd2362, -32'd7471, 32'd263},
{-32'd2266, 32'd820, 32'd1420, -32'd4217},
{-32'd6285, -32'd4600, 32'd771, -32'd13178},
{32'd4513, -32'd3710, -32'd4801, 32'd2971},
{32'd3000, 32'd2589, 32'd3248, -32'd4687},
{32'd7660, 32'd2643, -32'd507, -32'd3556},
{32'd10972, -32'd2010, 32'd9657, 32'd12485},
{-32'd3171, -32'd5326, -32'd5191, 32'd8927},
{-32'd540, 32'd2034, -32'd2461, -32'd5598},
{-32'd10403, 32'd2609, -32'd1620, 32'd1255},
{-32'd5415, -32'd2213, -32'd4851, -32'd3851},
{-32'd2577, 32'd10278, -32'd2819, -32'd3895},
{-32'd1843, 32'd13900, -32'd22412, -32'd7004},
{32'd2850, 32'd341, -32'd8946, -32'd7562},
{-32'd3148, 32'd3409, -32'd2647, 32'd292},
{32'd11200, 32'd3976, -32'd8463, -32'd2733},
{32'd4479, 32'd2717, 32'd8091, 32'd1179},
{32'd8760, 32'd12677, -32'd6254, 32'd5781},
{-32'd4256, 32'd1897, 32'd6569, 32'd6834},
{32'd12536, 32'd6369, -32'd3484, 32'd2119},
{32'd3577, -32'd46, -32'd5375, 32'd1518},
{32'd17804, 32'd8519, -32'd5928, 32'd2054},
{-32'd8613, -32'd5736, -32'd1254, -32'd4488},
{32'd10914, -32'd4070, 32'd355, 32'd5804},
{-32'd225, 32'd4342, -32'd2972, -32'd10658},
{32'd4358, 32'd6691, -32'd10355, 32'd631},
{-32'd4239, 32'd11249, 32'd1496, 32'd123},
{-32'd1865, -32'd3174, 32'd2130, -32'd1567},
{-32'd1556, 32'd8219, 32'd5092, -32'd2318},
{-32'd9638, 32'd3921, -32'd445, -32'd1588},
{-32'd410, 32'd9184, 32'd1919, -32'd1186},
{32'd2945, 32'd4924, -32'd1, -32'd5165},
{32'd13409, 32'd9325, -32'd10899, -32'd5496},
{32'd2346, 32'd10216, -32'd4514, -32'd1069},
{32'd103, -32'd8473, 32'd1244, 32'd6438},
{32'd2455, -32'd7519, 32'd15739, 32'd315},
{-32'd14322, -32'd9457, 32'd5544, 32'd1018},
{-32'd9853, 32'd2688, 32'd4515, 32'd1082},
{32'd9940, 32'd4935, 32'd7902, -32'd4422},
{-32'd1241, -32'd3563, -32'd6523, -32'd2498},
{-32'd5712, -32'd2004, -32'd1663, -32'd6325},
{-32'd6904, -32'd5876, 32'd10738, -32'd14955},
{32'd4817, -32'd5257, 32'd3411, 32'd5937},
{32'd323, 32'd5847, -32'd10542, -32'd8672},
{32'd4282, 32'd11714, -32'd8479, 32'd187},
{32'd4095, 32'd4824, 32'd14825, -32'd105},
{32'd9708, -32'd4963, -32'd1630, -32'd3299},
{-32'd2295, 32'd8100, -32'd3529, -32'd9552},
{32'd5404, 32'd961, 32'd5319, 32'd12426},
{32'd9622, 32'd6673, -32'd3483, -32'd1714},
{32'd3749, 32'd11127, 32'd78, 32'd1169},
{32'd3585, -32'd443, 32'd3280, -32'd4241},
{-32'd8985, -32'd2843, -32'd5027, -32'd8915},
{-32'd3907, -32'd3216, 32'd3681, -32'd1516},
{32'd12251, -32'd197, 32'd3992, -32'd764},
{32'd5535, 32'd4538, 32'd6950, -32'd1429},
{-32'd3553, -32'd1373, -32'd1305, 32'd1563},
{-32'd3384, 32'd4530, -32'd7291, 32'd7771},
{-32'd124, 32'd4033, 32'd6936, -32'd13614},
{32'd8170, -32'd15120, 32'd1820, -32'd1443},
{-32'd4493, 32'd3008, -32'd1618, -32'd2797},
{-32'd1984, 32'd4664, -32'd12163, -32'd7441},
{32'd6780, -32'd3183, -32'd3045, -32'd6586},
{32'd9544, 32'd11087, 32'd5499, -32'd9043},
{32'd753, 32'd2567, -32'd7223, 32'd6944},
{-32'd3523, 32'd10329, -32'd6530, 32'd1008},
{-32'd10591, 32'd3142, 32'd8971, 32'd5197},
{-32'd1013, 32'd8149, 32'd248, -32'd734},
{32'd3837, -32'd5378, 32'd1481, -32'd8866},
{32'd5662, 32'd5910, 32'd5165, -32'd71},
{32'd2276, 32'd8827, -32'd3322, 32'd867},
{32'd9758, 32'd10158, -32'd4259, 32'd5936},
{-32'd4069, -32'd569, -32'd7999, -32'd2969},
{32'd2851, 32'd186, -32'd9165, 32'd8143},
{32'd8971, -32'd3629, -32'd5164, -32'd5596},
{32'd13392, 32'd9010, 32'd1022, -32'd6857},
{-32'd3279, 32'd1033, -32'd3177, 32'd2587},
{32'd10478, 32'd26, -32'd3048, 32'd3396},
{-32'd10421, 32'd656, -32'd1597, 32'd14341},
{-32'd9963, 32'd4808, -32'd6871, -32'd1360},
{32'd2927, 32'd9650, -32'd676, -32'd139},
{-32'd3273, -32'd15485, -32'd852, 32'd1748},
{-32'd1638, -32'd7250, -32'd8828, -32'd1390},
{-32'd5299, -32'd6874, -32'd1859, 32'd9510},
{-32'd3677, 32'd6880, -32'd1821, -32'd6867},
{32'd4298, 32'd6849, 32'd2908, -32'd7009},
{32'd12384, 32'd3207, -32'd12028, 32'd8211},
{-32'd12335, 32'd835, -32'd18839, -32'd984},
{-32'd6563, 32'd14514, -32'd3121, 32'd6459},
{-32'd15216, -32'd1908, -32'd1706, -32'd3288},
{32'd10132, 32'd8636, 32'd11479, 32'd3590},
{-32'd4840, -32'd6368, -32'd1659, -32'd6502},
{32'd2245, 32'd3168, 32'd3107, -32'd7180},
{32'd16946, 32'd1279, 32'd2960, -32'd7822},
{-32'd3807, -32'd7600, -32'd5871, 32'd5433},
{-32'd4067, -32'd9698, 32'd2264, -32'd13289},
{32'd4227, 32'd14441, -32'd2458, -32'd911},
{32'd10457, 32'd3397, 32'd2782, -32'd248},
{-32'd1395, 32'd4364, -32'd1342, -32'd1628},
{-32'd3537, -32'd522, -32'd5821, -32'd10120},
{32'd16225, 32'd311, 32'd2211, -32'd3902},
{32'd8367, 32'd1129, -32'd2490, -32'd11395},
{-32'd16282, -32'd13530, 32'd1247, 32'd2494},
{-32'd97, 32'd1444, 32'd12298, 32'd12749},
{-32'd4213, -32'd6535, 32'd2724, 32'd11575},
{32'd3027, -32'd6051, 32'd6788, 32'd1327},
{-32'd15390, -32'd11135, -32'd3221, 32'd2002},
{32'd1388, -32'd10474, -32'd11397, 32'd6356},
{32'd5591, 32'd4539, 32'd2340, 32'd2835},
{32'd1252, -32'd5656, -32'd7289, 32'd4982},
{-32'd4751, 32'd2318, 32'd4528, 32'd213},
{-32'd1735, 32'd7660, 32'd1110, -32'd2569},
{-32'd9239, -32'd2040, -32'd20808, 32'd6287},
{32'd13453, 32'd10270, -32'd2025, -32'd6342},
{-32'd11928, 32'd6304, 32'd5435, 32'd7890},
{32'd3545, 32'd7311, -32'd6030, 32'd1890},
{32'd4769, -32'd1079, 32'd2461, -32'd5764},
{-32'd3716, -32'd6576, 32'd1182, -32'd11783},
{-32'd3155, -32'd4207, 32'd6787, -32'd10292},
{-32'd4875, -32'd604, -32'd11449, -32'd480},
{-32'd8091, -32'd6033, -32'd4049, 32'd6253},
{-32'd7046, -32'd1077, -32'd3339, -32'd3451},
{32'd3192, 32'd3689, 32'd9886, 32'd1997},
{32'd1707, -32'd1863, 32'd7583, 32'd7005},
{32'd13496, 32'd4039, 32'd7560, 32'd4003},
{-32'd3076, 32'd3397, -32'd2869, -32'd625},
{-32'd5628, 32'd9063, -32'd3107, 32'd1980},
{-32'd5078, -32'd8262, 32'd5479, -32'd2251},
{32'd14277, -32'd5770, 32'd2871, -32'd408},
{-32'd4694, -32'd4755, -32'd6880, -32'd1599},
{32'd1318, 32'd1075, -32'd6898, 32'd4246},
{-32'd16816, -32'd6556, -32'd7690, 32'd9175},
{32'd11081, -32'd6446, 32'd4101, -32'd6583},
{32'd2592, -32'd4455, 32'd842, 32'd9538},
{-32'd8559, -32'd8775, 32'd5305, 32'd9457},
{-32'd5003, 32'd10277, 32'd4524, 32'd9710},
{32'd122, -32'd9183, 32'd3159, 32'd1826},
{32'd5468, -32'd3013, 32'd3966, -32'd3226},
{32'd8802, 32'd188, 32'd3765, 32'd4885},
{32'd12091, -32'd721, -32'd4671, 32'd4911},
{32'd9016, 32'd6611, -32'd7437, -32'd4828},
{-32'd7104, -32'd10074, -32'd5978, 32'd6568},
{32'd4063, 32'd13425, -32'd965, -32'd1842},
{32'd1328, -32'd6080, -32'd6130, 32'd801},
{32'd9106, 32'd7564, -32'd2680, 32'd1611},
{32'd2482, 32'd20025, 32'd3348, -32'd3965},
{32'd3146, -32'd9892, 32'd3349, 32'd1586},
{-32'd6292, 32'd929, 32'd2759, 32'd6977},
{-32'd7269, -32'd5840, -32'd5937, -32'd2786},
{-32'd4415, -32'd4241, 32'd5624, 32'd2443},
{-32'd1657, 32'd2387, -32'd12465, 32'd5096},
{-32'd2088, -32'd5311, 32'd5403, 32'd4443},
{-32'd7074, -32'd6786, -32'd5085, 32'd88},
{32'd2488, 32'd416, -32'd6850, 32'd13075},
{32'd11160, -32'd486, 32'd6904, 32'd4155},
{32'd13811, 32'd4568, 32'd5886, 32'd10440},
{32'd1226, -32'd567, 32'd174, -32'd4413},
{-32'd7776, -32'd3278, 32'd4228, 32'd8636},
{32'd1919, 32'd5889, -32'd2025, 32'd15223},
{-32'd2360, -32'd4229, 32'd2102, -32'd225},
{32'd3850, -32'd3493, 32'd3672, 32'd4647},
{32'd3947, 32'd2685, 32'd1994, 32'd1823},
{32'd9240, 32'd9411, 32'd8686, -32'd4939},
{-32'd2219, -32'd4529, 32'd1815, -32'd6481},
{-32'd5270, 32'd14481, -32'd3161, 32'd8731},
{32'd1188, -32'd2077, -32'd7867, -32'd4699},
{-32'd16527, -32'd4941, 32'd11857, 32'd276},
{-32'd9102, -32'd8397, 32'd2292, -32'd3624},
{32'd3498, -32'd3565, 32'd6887, 32'd11747},
{32'd2789, 32'd2628, 32'd3473, -32'd4692},
{-32'd3673, -32'd1416, 32'd8138, 32'd13108},
{-32'd14184, -32'd179, -32'd382, 32'd2423},
{-32'd7622, -32'd10046, -32'd2775, 32'd9256},
{32'd1779, 32'd12848, -32'd2167, 32'd4258},
{32'd21884, 32'd4620, -32'd10446, 32'd6629},
{-32'd2419, -32'd6037, 32'd7264, 32'd6148},
{-32'd2501, 32'd9757, -32'd8106, -32'd5982},
{32'd5128, -32'd2180, -32'd3831, 32'd6454},
{32'd735, -32'd2417, 32'd2094, -32'd9230},
{32'd1401, 32'd6127, -32'd5994, -32'd9991},
{-32'd15112, -32'd7099, 32'd16720, 32'd1880},
{-32'd425, -32'd5594, 32'd4191, 32'd337},
{32'd4180, -32'd2136, 32'd4289, 32'd6379},
{32'd491, -32'd1116, 32'd2576, 32'd1910},
{32'd2962, 32'd2958, -32'd1593, -32'd3151},
{32'd3557, 32'd4192, -32'd8285, -32'd4799},
{-32'd4897, 32'd134, 32'd3146, 32'd1621},
{32'd624, -32'd1470, -32'd9066, -32'd11852},
{32'd1155, -32'd9200, 32'd6500, -32'd7644},
{-32'd957, -32'd4120, 32'd9203, -32'd112},
{32'd1270, -32'd3651, -32'd5203, 32'd5966},
{32'd4770, 32'd357, -32'd619, 32'd611},
{-32'd1667, 32'd12492, -32'd10134, 32'd822},
{-32'd11943, 32'd2602, -32'd3813, 32'd6704},
{-32'd3073, -32'd917, -32'd4654, -32'd7796},
{32'd3238, -32'd2754, 32'd3167, -32'd5367},
{32'd6044, 32'd3843, -32'd920, 32'd5099},
{-32'd176, 32'd6054, -32'd6856, 32'd4203},
{32'd6219, 32'd6822, 32'd7060, 32'd9265},
{32'd749, 32'd4793, 32'd7624, -32'd8710},
{-32'd4834, 32'd859, 32'd4109, -32'd2567},
{-32'd8493, -32'd2718, 32'd1544, -32'd14159},
{32'd6124, 32'd696, -32'd10421, 32'd7191},
{32'd2642, 32'd6707, 32'd3784, -32'd3370},
{-32'd2665, -32'd9328, 32'd22545, 32'd10795},
{-32'd1521, -32'd1175, -32'd6406, 32'd5827},
{-32'd1675, -32'd5928, 32'd4017, 32'd7140},
{-32'd535, 32'd4986, 32'd1034, -32'd3905},
{32'd7882, 32'd4551, 32'd10548, -32'd2706},
{32'd5879, 32'd373, 32'd8038, -32'd3366},
{-32'd10192, -32'd7223, -32'd6417, 32'd3369},
{32'd1570, -32'd711, 32'd14517, -32'd2988},
{32'd13158, -32'd2369, 32'd11920, 32'd7992},
{32'd3435, -32'd3101, 32'd2451, 32'd3101},
{32'd18132, -32'd534, 32'd3960, -32'd17191},
{-32'd9967, 32'd811, -32'd10223, -32'd2707},
{32'd14809, -32'd4350, 32'd3017, -32'd2241},
{-32'd5720, -32'd911, -32'd12561, -32'd2158},
{-32'd2450, 32'd288, 32'd1855, 32'd6225},
{-32'd10663, -32'd3065, 32'd2948, 32'd5335},
{32'd3025, -32'd9840, 32'd1625, -32'd3513},
{32'd13493, 32'd4831, -32'd858, -32'd6056},
{-32'd3585, 32'd7505, -32'd2648, 32'd4247},
{32'd17, 32'd2698, 32'd5557, 32'd4495},
{32'd1862, -32'd369, -32'd3602, -32'd8048},
{32'd3208, -32'd1648, 32'd6964, 32'd2470},
{32'd5923, -32'd8772, -32'd1582, -32'd2383},
{32'd2950, 32'd4222, 32'd2798, 32'd2967},
{32'd9271, 32'd5749, 32'd2635, 32'd433},
{32'd14746, 32'd38, 32'd83, 32'd863},
{-32'd4948, 32'd2867, -32'd3529, -32'd3218},
{32'd3251, -32'd5262, 32'd2508, -32'd18398},
{32'd15626, 32'd12196, -32'd10490, 32'd876},
{32'd2075, -32'd743, -32'd9316, -32'd5764},
{32'd2346, 32'd4093, -32'd1133, 32'd1988},
{32'd6901, 32'd9544, -32'd10480, 32'd1744},
{32'd1847, 32'd1747, -32'd748, -32'd596},
{32'd4655, -32'd11117, 32'd905, -32'd4572},
{32'd2000, 32'd725, 32'd2946, -32'd1125},
{32'd4456, 32'd4432, 32'd7963, 32'd636},
{-32'd4881, 32'd6392, 32'd3838, -32'd5693},
{-32'd5846, 32'd5739, -32'd4637, 32'd200},
{32'd1618, -32'd1034, -32'd3140, -32'd4364},
{-32'd1698, 32'd8735, 32'd1691, 32'd3388},
{-32'd906, -32'd6068, 32'd6219, -32'd13762},
{-32'd6943, -32'd7933, 32'd1741, -32'd1961},
{-32'd11450, -32'd10719, -32'd9615, -32'd3417},
{-32'd4598, -32'd4796, 32'd1971, 32'd7261},
{32'd4323, -32'd12230, -32'd5638, -32'd4017},
{32'd4812, 32'd3111, 32'd8129, 32'd7209},
{32'd7921, -32'd6934, 32'd5932, 32'd694},
{32'd7542, 32'd2357, -32'd3486, 32'd1660}
},
{{32'd3545, -32'd2867, -32'd3002, -32'd3602},
{-32'd5600, -32'd4969, 32'd212, 32'd10499},
{-32'd11660, 32'd3902, 32'd7111, -32'd105},
{-32'd1878, -32'd3836, 32'd1913, 32'd7225},
{32'd5376, 32'd8397, 32'd2571, 32'd1020},
{-32'd4624, 32'd2635, -32'd2234, 32'd984},
{-32'd7392, -32'd4991, -32'd3159, 32'd4185},
{32'd2316, -32'd4955, -32'd1166, -32'd749},
{-32'd2136, -32'd3702, 32'd16, 32'd8336},
{32'd13537, 32'd8873, 32'd3900, 32'd2334},
{32'd2195, 32'd1258, 32'd3584, 32'd4327},
{32'd2916, -32'd32, 32'd719, -32'd4660},
{-32'd4944, -32'd9429, -32'd8618, -32'd2700},
{32'd2894, -32'd6589, -32'd2446, -32'd303},
{32'd6761, -32'd9132, -32'd1391, -32'd2602},
{32'd10849, 32'd355, -32'd882, -32'd17000},
{32'd2035, 32'd1248, 32'd7074, -32'd2711},
{32'd958, 32'd4239, -32'd7423, 32'd8946},
{32'd9339, 32'd1582, 32'd5006, -32'd9114},
{32'd2126, 32'd674, 32'd11694, -32'd8957},
{-32'd2235, 32'd1788, 32'd4258, 32'd3277},
{-32'd11479, -32'd8040, 32'd3399, -32'd3182},
{-32'd10218, -32'd4116, 32'd1532, -32'd233},
{-32'd3891, -32'd1997, -32'd3478, -32'd566},
{32'd6722, 32'd2591, 32'd5834, 32'd1518},
{-32'd12484, -32'd8897, 32'd88, -32'd772},
{32'd4768, -32'd7443, 32'd2313, 32'd2216},
{32'd6058, 32'd8273, -32'd2576, -32'd21},
{-32'd2909, 32'd10796, 32'd1016, -32'd7330},
{-32'd5148, 32'd3060, -32'd6358, -32'd1663},
{-32'd1299, 32'd1481, 32'd883, -32'd471},
{-32'd6877, 32'd708, -32'd3148, 32'd4277},
{32'd2772, 32'd6191, 32'd3534, -32'd3699},
{32'd466, -32'd3512, -32'd2494, -32'd1846},
{32'd5292, 32'd5880, 32'd3318, 32'd98},
{32'd5002, -32'd7171, 32'd3818, 32'd1803},
{-32'd6224, -32'd2893, -32'd9855, 32'd6906},
{-32'd9656, -32'd5529, 32'd687, -32'd12627},
{-32'd438, 32'd5606, -32'd2607, 32'd2433},
{32'd10515, 32'd11038, 32'd2344, 32'd518},
{-32'd842, -32'd12709, -32'd701, -32'd4622},
{32'd13181, 32'd350, -32'd3961, 32'd2996},
{32'd14668, -32'd485, 32'd8580, -32'd13266},
{-32'd1136, 32'd2173, -32'd3511, -32'd1655},
{-32'd5770, -32'd11682, -32'd3760, -32'd8972},
{32'd6965, -32'd303, -32'd5205, -32'd7622},
{-32'd7892, -32'd3860, 32'd6306, -32'd5976},
{-32'd2088, 32'd1449, -32'd758, 32'd171},
{32'd413, 32'd2260, 32'd3862, 32'd3766},
{-32'd2490, 32'd5274, -32'd4745, -32'd11001},
{-32'd7125, -32'd12035, 32'd2907, 32'd5135},
{32'd1064, 32'd5113, -32'd7617, 32'd5263},
{-32'd5452, 32'd1014, -32'd1968, -32'd1533},
{-32'd7230, -32'd2227, 32'd10610, 32'd3067},
{-32'd5564, 32'd1298, -32'd9579, -32'd8007},
{-32'd10230, -32'd1958, -32'd1357, -32'd747},
{32'd2237, 32'd9850, 32'd8741, 32'd6691},
{-32'd5482, -32'd3330, 32'd2944, -32'd8435},
{32'd1283, 32'd6, 32'd4603, -32'd1856},
{32'd6212, 32'd6538, 32'd782, 32'd2235},
{32'd923, -32'd900, -32'd1721, 32'd7872},
{-32'd755, -32'd7731, -32'd7803, -32'd10182},
{32'd3564, -32'd4003, -32'd575, -32'd1246},
{32'd7, -32'd5133, 32'd2634, 32'd4147},
{32'd680, 32'd771, -32'd4172, 32'd3589},
{-32'd3159, 32'd7816, -32'd1891, 32'd5952},
{-32'd1166, -32'd6462, 32'd2957, -32'd11945},
{-32'd13508, 32'd6619, -32'd6230, 32'd6442},
{32'd11279, 32'd16395, -32'd11891, -32'd3371},
{-32'd1888, -32'd3935, -32'd5324, 32'd7192},
{-32'd479, 32'd12254, -32'd9962, -32'd3260},
{32'd3450, 32'd10546, -32'd10185, -32'd3398},
{-32'd7305, 32'd1696, -32'd12229, 32'd8615},
{-32'd5398, 32'd3914, -32'd6556, -32'd6410},
{32'd3286, 32'd2435, 32'd1928, -32'd793},
{-32'd1315, -32'd10216, -32'd755, -32'd4223},
{-32'd569, -32'd12659, 32'd4273, -32'd9468},
{32'd13957, 32'd5200, -32'd2846, -32'd10052},
{32'd8389, 32'd5832, -32'd6912, 32'd10862},
{-32'd1449, 32'd2162, 32'd5808, 32'd11624},
{32'd4524, 32'd15035, -32'd83, 32'd4675},
{32'd5771, 32'd5980, 32'd4811, 32'd6622},
{-32'd5039, -32'd2804, 32'd8616, -32'd1083},
{-32'd2139, -32'd3926, 32'd1950, -32'd6866},
{-32'd11114, 32'd4660, 32'd2661, 32'd5339},
{-32'd7359, 32'd5705, -32'd3550, -32'd13814},
{-32'd3371, -32'd3340, -32'd975, -32'd4554},
{-32'd4503, -32'd13327, -32'd2476, 32'd6705},
{32'd13265, -32'd7287, 32'd7876, -32'd3947},
{-32'd7518, -32'd4871, 32'd7347, 32'd464},
{32'd5504, 32'd11288, 32'd2431, 32'd5488},
{32'd20, -32'd4036, -32'd11562, 32'd1730},
{32'd6410, 32'd9929, -32'd3410, 32'd1936},
{32'd1250, 32'd5993, 32'd2383, 32'd8356},
{-32'd2857, -32'd3502, -32'd2343, 32'd5783},
{-32'd324, 32'd7253, -32'd9922, 32'd3181},
{32'd16734, 32'd14609, 32'd1417, -32'd1198},
{-32'd10320, 32'd3513, 32'd1575, -32'd1041},
{-32'd18188, 32'd1746, -32'd6602, 32'd7835},
{32'd3522, 32'd13792, 32'd6534, -32'd3009},
{-32'd9825, -32'd2168, -32'd5845, -32'd14952},
{-32'd4802, 32'd44, -32'd7129, -32'd2163},
{32'd1457, -32'd11518, 32'd9058, -32'd2355},
{32'd5364, 32'd4822, 32'd1492, -32'd9704},
{32'd10658, 32'd6538, 32'd6094, -32'd3006},
{32'd5432, 32'd3503, -32'd5345, -32'd783},
{-32'd977, 32'd2847, 32'd7064, -32'd8660},
{-32'd8860, 32'd378, 32'd865, -32'd2096},
{32'd9496, -32'd1074, 32'd2192, -32'd6365},
{32'd12407, 32'd79, -32'd3403, -32'd4845},
{32'd4348, -32'd3033, -32'd2615, 32'd3036},
{32'd1816, 32'd6681, 32'd14345, -32'd403},
{32'd3278, 32'd3158, 32'd8352, 32'd3495},
{32'd15135, 32'd13556, 32'd9813, -32'd1335},
{-32'd6210, -32'd13142, 32'd1294, -32'd3841},
{32'd3756, -32'd7696, -32'd10159, 32'd68},
{32'd1163, 32'd2655, 32'd9323, -32'd5098},
{32'd3465, 32'd8760, 32'd273, -32'd5554},
{32'd13814, 32'd10786, 32'd3498, -32'd81},
{32'd9185, 32'd12122, 32'd3940, 32'd1272},
{32'd2264, -32'd5903, -32'd2633, 32'd3433},
{-32'd1191, 32'd203, 32'd8448, -32'd3778},
{-32'd2038, 32'd9246, -32'd8316, -32'd6900},
{-32'd3903, -32'd499, 32'd3967, -32'd2461},
{-32'd4584, 32'd9070, 32'd5496, 32'd7871},
{-32'd6890, -32'd444, -32'd4998, 32'd7264},
{32'd8884, -32'd8094, 32'd1145, 32'd7744},
{-32'd1203, 32'd2077, -32'd1988, 32'd4838},
{-32'd9379, -32'd3866, -32'd358, 32'd6738},
{-32'd5669, 32'd1149, -32'd7282, 32'd3961},
{32'd4247, -32'd5799, -32'd3306, -32'd10858},
{-32'd4505, -32'd1899, -32'd10764, -32'd4989},
{-32'd827, -32'd13390, -32'd12601, -32'd5804},
{-32'd10730, 32'd7994, -32'd3729, 32'd11124},
{32'd198, 32'd2499, -32'd111, 32'd4025},
{32'd10256, 32'd11814, -32'd2136, 32'd957},
{32'd7417, -32'd1808, -32'd634, 32'd1649},
{-32'd7779, -32'd2235, 32'd2324, -32'd5677},
{32'd6545, 32'd3640, 32'd12334, -32'd1570},
{-32'd8710, -32'd10131, -32'd9649, -32'd4348},
{32'd4949, 32'd5906, 32'd8381, -32'd3503},
{-32'd2187, 32'd2448, 32'd8576, 32'd1628},
{32'd110, 32'd779, -32'd15018, 32'd5001},
{-32'd16190, 32'd726, -32'd4225, -32'd5441},
{32'd1717, 32'd1592, 32'd1061, 32'd8359},
{32'd9194, 32'd11418, -32'd5879, 32'd5412},
{-32'd7371, 32'd3878, 32'd3780, 32'd2064},
{-32'd2949, 32'd8746, -32'd774, 32'd2835},
{-32'd4302, -32'd2103, 32'd1814, 32'd6330},
{-32'd5778, 32'd3316, 32'd688, 32'd3377},
{-32'd1498, -32'd2776, 32'd1298, -32'd7311},
{32'd3776, 32'd4570, 32'd8119, -32'd14429},
{32'd3750, 32'd788, -32'd6660, -32'd8970},
{32'd2268, -32'd3413, 32'd7672, -32'd3229},
{-32'd10755, -32'd8070, 32'd2932, -32'd5859},
{-32'd8242, -32'd6736, 32'd3876, 32'd3653},
{32'd9671, 32'd7695, 32'd2358, -32'd2041},
{-32'd9301, -32'd8079, 32'd5118, 32'd1165},
{-32'd14472, 32'd841, -32'd2740, -32'd5254},
{32'd17157, 32'd11592, -32'd22, -32'd9403},
{32'd4094, -32'd1135, -32'd3504, -32'd2236},
{32'd2201, 32'd5062, 32'd9568, -32'd9243},
{-32'd8028, 32'd3453, 32'd2249, -32'd9914},
{-32'd1731, 32'd2700, 32'd2867, 32'd2503},
{32'd1964, 32'd5021, -32'd12391, -32'd2154},
{-32'd2727, -32'd12854, -32'd6032, -32'd4157},
{-32'd4133, -32'd6899, 32'd2014, -32'd6996},
{32'd2959, -32'd9386, -32'd5799, 32'd3697},
{-32'd12270, 32'd256, -32'd1651, 32'd3360},
{-32'd4527, 32'd6156, -32'd1078, 32'd1962},
{32'd3422, -32'd3242, 32'd2619, 32'd6041},
{-32'd10122, -32'd333, 32'd7105, 32'd7808},
{32'd4827, 32'd4524, 32'd725, 32'd2985},
{-32'd5252, -32'd3975, -32'd3520, 32'd2993},
{-32'd3211, 32'd10735, 32'd8708, 32'd6429},
{-32'd8449, -32'd602, -32'd1973, -32'd9602},
{32'd11599, -32'd6874, 32'd6981, 32'd10546},
{-32'd2133, 32'd7618, 32'd1735, -32'd1895},
{32'd9258, 32'd1510, 32'd8313, 32'd2730},
{-32'd10018, -32'd4664, 32'd1712, -32'd348},
{32'd5259, 32'd6888, -32'd6848, -32'd7450},
{-32'd1442, -32'd254, -32'd8812, -32'd2005},
{-32'd2843, 32'd4853, -32'd5312, -32'd10339},
{32'd3881, 32'd1504, 32'd97, -32'd8168},
{-32'd4144, 32'd1131, 32'd7144, 32'd3850},
{-32'd5092, 32'd991, 32'd4716, 32'd12455},
{32'd4459, -32'd259, -32'd4697, 32'd4370},
{-32'd14795, 32'd7178, -32'd6478, 32'd3907},
{32'd113, 32'd664, -32'd1683, 32'd12127},
{32'd958, 32'd2395, -32'd550, -32'd5773},
{-32'd9034, -32'd3053, 32'd1157, -32'd1275},
{-32'd3930, -32'd3076, -32'd7188, 32'd2868},
{32'd195, -32'd4992, -32'd7461, 32'd8822},
{-32'd7259, -32'd3661, 32'd3527, 32'd11250},
{32'd7886, 32'd3404, -32'd8637, 32'd491},
{32'd129, 32'd2907, 32'd4958, 32'd5033},
{-32'd4076, 32'd914, 32'd8168, 32'd9518},
{-32'd1718, 32'd4704, -32'd7333, -32'd4601},
{-32'd8007, 32'd5159, -32'd4850, 32'd6148},
{-32'd3008, -32'd5119, -32'd223, -32'd3084},
{-32'd5848, -32'd5697, -32'd335, -32'd6787},
{32'd6651, 32'd7741, -32'd1013, -32'd6242},
{32'd3959, 32'd777, 32'd4094, -32'd1284},
{32'd289, -32'd5656, 32'd5645, 32'd9584},
{-32'd11721, -32'd4925, 32'd2244, -32'd5883},
{-32'd3762, 32'd13286, 32'd3650, -32'd154},
{32'd4913, -32'd4210, -32'd251, -32'd6972},
{-32'd8507, 32'd1261, 32'd448, 32'd4581},
{32'd5897, 32'd4968, 32'd10481, 32'd6738},
{32'd4914, 32'd2205, 32'd2570, -32'd5375},
{-32'd1062, -32'd4947, -32'd8197, -32'd45},
{32'd6142, -32'd3036, -32'd3587, -32'd2154},
{-32'd12811, 32'd4087, -32'd7959, -32'd10812},
{32'd1970, 32'd4408, -32'd368, -32'd1407},
{-32'd2301, -32'd8533, 32'd6734, -32'd8237},
{-32'd44, -32'd4100, 32'd3798, -32'd337},
{32'd4232, 32'd5914, -32'd3943, 32'd12985},
{-32'd19002, -32'd6194, -32'd12116, 32'd56},
{32'd12166, 32'd13548, 32'd1234, -32'd4965},
{-32'd8596, 32'd2360, 32'd6002, -32'd5610},
{32'd10043, 32'd2383, -32'd744, -32'd6937},
{32'd5297, 32'd427, 32'd6216, -32'd1654},
{32'd10608, 32'd7541, 32'd8825, 32'd2306},
{32'd671, 32'd6320, 32'd4190, 32'd5423},
{32'd4787, -32'd756, -32'd1120, 32'd1337},
{-32'd503, 32'd8808, 32'd3265, 32'd723},
{32'd11411, -32'd1736, 32'd8242, -32'd11023},
{-32'd4377, -32'd5965, -32'd1436, 32'd10538},
{32'd14115, 32'd1138, -32'd705, -32'd2896},
{-32'd5451, -32'd8208, 32'd1557, 32'd86},
{-32'd2225, 32'd3388, 32'd1703, -32'd1172},
{-32'd7917, -32'd1522, -32'd3956, 32'd6068},
{-32'd8435, 32'd6091, -32'd2448, -32'd600},
{32'd4500, -32'd13970, -32'd6683, 32'd3246},
{-32'd11085, -32'd2792, 32'd1045, 32'd4982},
{-32'd11360, -32'd10087, -32'd4702, -32'd128},
{32'd1944, -32'd964, 32'd1212, 32'd1575},
{-32'd10581, 32'd3154, -32'd8809, 32'd841},
{32'd8380, 32'd5248, -32'd1592, 32'd1031},
{-32'd6805, -32'd2351, -32'd7731, -32'd5750},
{32'd68, -32'd2199, 32'd2339, -32'd2057},
{32'd3150, -32'd2863, -32'd5178, -32'd13778},
{-32'd7384, -32'd14230, -32'd459, 32'd356},
{-32'd2814, -32'd1134, -32'd395, 32'd2564},
{32'd9007, 32'd4205, 32'd2816, 32'd2009},
{32'd456, -32'd9739, 32'd2398, 32'd14163},
{-32'd3391, -32'd1047, 32'd1452, -32'd3614},
{32'd5404, 32'd3637, 32'd5983, -32'd1100},
{-32'd373, 32'd4076, 32'd3104, -32'd6557},
{-32'd3649, -32'd6171, -32'd1638, -32'd803},
{-32'd4492, -32'd3123, -32'd3642, 32'd1095},
{-32'd4018, 32'd7203, 32'd6023, -32'd1040},
{32'd1006, 32'd2107, -32'd3978, 32'd1684},
{32'd2908, -32'd479, 32'd4088, 32'd6869},
{-32'd4429, -32'd5665, 32'd3262, -32'd17018},
{-32'd883, -32'd4365, 32'd14599, 32'd3764},
{-32'd3644, -32'd5092, 32'd11751, 32'd3313},
{-32'd1793, 32'd10387, 32'd484, -32'd723},
{-32'd14720, -32'd3550, -32'd2042, -32'd6536},
{32'd4209, 32'd2098, 32'd4020, -32'd434},
{-32'd13164, 32'd37, 32'd2133, 32'd12545},
{32'd2462, 32'd2128, -32'd3267, 32'd7426},
{-32'd9340, -32'd1872, 32'd7204, -32'd8620},
{32'd4902, 32'd871, 32'd1512, -32'd9676},
{-32'd12049, -32'd713, 32'd5399, 32'd11523},
{-32'd3256, 32'd3872, 32'd220, -32'd7814},
{32'd12187, 32'd6752, 32'd155, 32'd7831},
{-32'd438, -32'd4985, -32'd2228, 32'd1920},
{-32'd7591, -32'd10162, 32'd778, -32'd6208},
{-32'd9006, 32'd813, 32'd850, 32'd3823},
{-32'd423, 32'd11253, -32'd5116, -32'd2967},
{-32'd17266, 32'd4874, -32'd4918, 32'd7192},
{-32'd6796, 32'd11182, 32'd3551, -32'd4283},
{-32'd5654, -32'd6593, -32'd12034, -32'd847},
{-32'd2382, -32'd2076, -32'd5767, -32'd11010},
{32'd10853, -32'd8536, 32'd2093, 32'd2515},
{32'd8742, 32'd8362, 32'd1534, 32'd5754},
{32'd10626, 32'd8957, -32'd15798, -32'd5095},
{-32'd4991, -32'd11757, -32'd7225, -32'd8544},
{-32'd1911, 32'd2417, -32'd5255, -32'd8782},
{-32'd1664, 32'd14387, 32'd13614, 32'd3489},
{32'd13674, 32'd2400, -32'd4978, 32'd4272},
{32'd10781, 32'd9913, -32'd3041, 32'd7885},
{-32'd2559, 32'd4557, -32'd9193, 32'd6703},
{-32'd1056, -32'd952, -32'd3519, 32'd9363},
{-32'd914, -32'd3761, 32'd5548, -32'd9174},
{-32'd309, -32'd720, 32'd4162, 32'd3326},
{-32'd12078, -32'd3264, 32'd5966, -32'd9903},
{32'd7543, -32'd1488, -32'd7382, -32'd2958},
{-32'd2089, 32'd3276, 32'd1920, -32'd414},
{-32'd4363, -32'd11397, -32'd1120, 32'd949},
{32'd5094, 32'd1314, 32'd398, 32'd7866},
{-32'd1957, 32'd5375, 32'd4735, -32'd12764},
{-32'd4757, -32'd12362, -32'd7506, -32'd7005},
{-32'd10192, -32'd3199, -32'd9861, 32'd1032},
{-32'd5169, -32'd2945, -32'd358, -32'd3826},
{32'd182, -32'd9844, 32'd3219, 32'd1594},
{32'd5321, 32'd4098, -32'd3542, -32'd9434},
{32'd5604, 32'd5180, 32'd3785, 32'd3749},
{32'd8170, -32'd5553, -32'd5721, -32'd8361}
},
{{-32'd10728, -32'd2903, 32'd6609, -32'd6270},
{32'd11502, -32'd6325, -32'd5509, -32'd4519},
{32'd7112, -32'd2725, 32'd14149, -32'd17418},
{32'd1861, -32'd18967, 32'd9491, -32'd9216},
{32'd3500, 32'd128, 32'd8510, 32'd3059},
{32'd2258, -32'd8175, 32'd4814, 32'd6225},
{32'd5762, -32'd5850, -32'd4623, 32'd1146},
{32'd6183, 32'd3015, 32'd4569, -32'd18036},
{32'd7411, 32'd5869, 32'd339, 32'd8464},
{32'd1279, 32'd1484, 32'd1686, -32'd1018},
{-32'd1383, -32'd9109, 32'd292, -32'd464},
{32'd12694, -32'd4399, -32'd2587, 32'd11741},
{-32'd17667, -32'd7952, -32'd1374, 32'd2942},
{-32'd1109, 32'd6078, -32'd9178, 32'd600},
{-32'd7137, -32'd7136, 32'd6650, 32'd659},
{-32'd6826, -32'd20855, 32'd254, 32'd13086},
{32'd9474, 32'd5945, 32'd609, -32'd11606},
{32'd14109, -32'd8874, 32'd15184, -32'd10066},
{-32'd12863, -32'd9101, 32'd7252, 32'd449},
{32'd1773, -32'd5893, -32'd6324, -32'd6517},
{-32'd5104, 32'd565, -32'd2005, -32'd8725},
{-32'd4839, -32'd5332, -32'd249, 32'd13652},
{-32'd6511, 32'd835, 32'd914, 32'd9851},
{-32'd8279, 32'd9705, -32'd6196, 32'd3071},
{32'd8119, 32'd5098, -32'd3724, -32'd1928},
{32'd1921, 32'd164, 32'd5062, -32'd17983},
{-32'd9864, -32'd1361, -32'd3281, 32'd9186},
{32'd4157, 32'd17546, 32'd8984, -32'd5278},
{32'd11709, 32'd17189, 32'd2090, -32'd27},
{-32'd9030, 32'd6783, 32'd12054, 32'd20783},
{32'd1618, -32'd2319, 32'd19154, -32'd15352},
{-32'd3942, 32'd3185, -32'd4229, 32'd975},
{-32'd1016, -32'd1219, -32'd6141, -32'd1961},
{-32'd4865, -32'd6996, -32'd287, 32'd5675},
{32'd8137, 32'd5796, 32'd6916, -32'd2921},
{-32'd8425, -32'd12281, -32'd6166, 32'd2779},
{32'd7685, 32'd4457, 32'd6623, -32'd25625},
{-32'd103, -32'd16735, 32'd1771, 32'd9113},
{32'd16738, 32'd14276, -32'd3052, -32'd6354},
{32'd14400, 32'd2301, -32'd4893, 32'd12197},
{32'd6589, -32'd8289, -32'd11278, 32'd2582},
{32'd5526, 32'd2650, -32'd13279, -32'd1892},
{-32'd5244, -32'd2040, 32'd4735, 32'd5507},
{-32'd17164, -32'd1527, 32'd6339, 32'd6018},
{-32'd20925, 32'd8695, 32'd5340, 32'd2321},
{32'd105, 32'd2560, -32'd2790, 32'd4826},
{-32'd2793, -32'd10491, 32'd729, 32'd6483},
{-32'd13613, -32'd9181, 32'd3056, 32'd3107},
{32'd516, 32'd6702, -32'd9280, 32'd2284},
{32'd9589, -32'd4943, -32'd12330, -32'd2433},
{32'd2248, 32'd5519, -32'd14625, -32'd8178},
{-32'd5071, 32'd5340, -32'd14526, -32'd6988},
{-32'd6244, -32'd6444, -32'd3716, 32'd8917},
{32'd5824, 32'd4947, -32'd9184, 32'd10568},
{-32'd2179, 32'd9261, 32'd8126, 32'd23020},
{32'd19041, 32'd13301, 32'd2366, -32'd20600},
{32'd20423, 32'd4356, 32'd6322, -32'd10464},
{32'd309, -32'd10749, -32'd4914, 32'd431},
{-32'd466, -32'd14247, 32'd990, 32'd6042},
{32'd12123, 32'd9844, 32'd10473, -32'd6933},
{32'd1157, -32'd112, -32'd1022, -32'd3158},
{32'd12978, 32'd9159, 32'd10375, 32'd3024},
{32'd1501, 32'd983, -32'd3062, -32'd1215},
{-32'd2239, 32'd4657, 32'd3209, -32'd588},
{-32'd10001, -32'd3509, -32'd8125, 32'd5741},
{32'd6719, 32'd2709, 32'd4065, 32'd604},
{-32'd12673, -32'd8353, -32'd4646, 32'd5022},
{32'd14611, 32'd4508, 32'd13649, -32'd2322},
{-32'd13577, -32'd11667, -32'd4758, -32'd4577},
{32'd12581, 32'd5471, -32'd592, -32'd2116},
{-32'd2871, 32'd2681, -32'd6627, -32'd8644},
{-32'd9823, -32'd5654, 32'd9001, -32'd9738},
{32'd121, 32'd13757, -32'd11156, -32'd2411},
{32'd1719, -32'd11432, -32'd1928, 32'd12566},
{32'd2292, 32'd17742, -32'd4159, 32'd2571},
{32'd613, 32'd17465, -32'd168, -32'd11437},
{32'd7985, 32'd558, 32'd13431, -32'd6189},
{32'd6138, -32'd2770, 32'd2203, 32'd4491},
{-32'd6743, 32'd11584, 32'd3825, -32'd4005},
{32'd2661, 32'd5720, 32'd2779, -32'd11354},
{32'd1204, -32'd2035, -32'd1788, -32'd4322},
{32'd2707, -32'd1474, 32'd7869, 32'd1178},
{32'd11938, -32'd5042, -32'd9407, 32'd5504},
{32'd10662, 32'd15634, -32'd8067, -32'd5621},
{-32'd4188, -32'd1636, 32'd3435, 32'd6662},
{-32'd1551, 32'd9920, 32'd989, -32'd4989},
{32'd4870, 32'd13119, 32'd5380, -32'd12749},
{-32'd6046, 32'd2442, -32'd1074, 32'd3652},
{-32'd2662, 32'd5553, 32'd382, -32'd12967},
{32'd812, 32'd10372, 32'd2136, -32'd2024},
{32'd5659, 32'd6234, -32'd35, 32'd7746},
{32'd4010, -32'd4692, -32'd10809, 32'd15473},
{-32'd2421, 32'd2536, 32'd7114, -32'd4053},
{32'd4357, -32'd13775, -32'd6002, -32'd8590},
{32'd8733, 32'd8778, 32'd11692, -32'd2902},
{-32'd2100, -32'd4453, 32'd11038, -32'd14993},
{32'd8382, -32'd2704, 32'd5367, -32'd1476},
{-32'd5891, -32'd7208, 32'd17356, 32'd2971},
{32'd4222, 32'd9305, -32'd3544, -32'd6460},
{-32'd4569, 32'd826, 32'd14031, 32'd6295},
{-32'd8536, -32'd7692, 32'd10334, -32'd7725},
{-32'd9908, 32'd8382, -32'd4605, 32'd11411},
{32'd7758, 32'd12180, 32'd9208, -32'd1968},
{-32'd12303, 32'd14264, -32'd1337, 32'd624},
{32'd6268, -32'd4522, -32'd6636, -32'd5017},
{32'd5023, -32'd15490, -32'd1570, 32'd3251},
{32'd788, 32'd12990, 32'd556, 32'd3311},
{-32'd8215, -32'd3117, -32'd6251, 32'd9371},
{-32'd14171, -32'd10160, 32'd584, 32'd5373},
{-32'd12479, -32'd16213, 32'd4326, -32'd5296},
{32'd12880, 32'd9582, -32'd5761, -32'd6161},
{32'd57, 32'd20960, 32'd1006, 32'd57},
{-32'd3464, -32'd8506, -32'd6379, -32'd178},
{-32'd1830, -32'd3543, 32'd14629, -32'd1475},
{32'd2757, -32'd13190, -32'd13779, 32'd12193},
{32'd7631, 32'd7479, 32'd1635, 32'd1953},
{32'd1103, 32'd12666, -32'd15633, -32'd4508},
{32'd9781, -32'd2641, 32'd4044, 32'd3595},
{-32'd7299, -32'd1900, -32'd1046, 32'd114},
{32'd10148, -32'd6471, -32'd717, -32'd5924},
{-32'd8386, -32'd9796, -32'd12686, 32'd5732},
{32'd1236, 32'd5672, -32'd8380, -32'd2672},
{32'd5748, -32'd5265, -32'd6597, -32'd1849},
{32'd12073, -32'd9751, 32'd21872, -32'd12392},
{-32'd7601, -32'd15374, 32'd8114, 32'd2213},
{32'd4385, 32'd24381, -32'd779, -32'd9153},
{-32'd6382, -32'd4024, 32'd1554, 32'd16764},
{32'd7824, 32'd9979, 32'd269, -32'd11456},
{-32'd2423, 32'd308, -32'd4437, 32'd11442},
{32'd2643, 32'd675, 32'd4849, -32'd15230},
{-32'd4376, 32'd2661, 32'd7865, 32'd5254},
{-32'd906, 32'd7761, 32'd3876, 32'd2353},
{-32'd1750, 32'd7654, 32'd10287, -32'd7704},
{32'd7327, 32'd6753, -32'd10630, -32'd908},
{-32'd1142, -32'd11212, -32'd15228, 32'd164},
{-32'd7211, -32'd4304, -32'd8326, -32'd1695},
{-32'd75, -32'd268, 32'd9530, -32'd8726},
{32'd6019, -32'd7151, -32'd548, -32'd9823},
{32'd12870, 32'd2473, 32'd9378, 32'd6365},
{-32'd8196, 32'd453, -32'd478, 32'd726},
{32'd6398, -32'd4862, -32'd9587, -32'd10033},
{-32'd3291, 32'd6420, 32'd13684, -32'd7755},
{32'd5153, 32'd344, -32'd12245, -32'd5328},
{-32'd2051, 32'd6782, -32'd6792, 32'd6564},
{32'd10932, 32'd15066, 32'd908, -32'd10988},
{32'd15230, 32'd9290, -32'd14275, -32'd526},
{32'd5163, -32'd6039, 32'd1033, -32'd1324},
{32'd11740, -32'd11499, -32'd5581, -32'd4505},
{32'd903, -32'd2896, 32'd4737, -32'd2056},
{-32'd3275, -32'd4659, 32'd7318, -32'd603},
{-32'd12983, 32'd6745, -32'd7173, 32'd318},
{-32'd10828, -32'd8169, -32'd18596, -32'd4686},
{32'd535, -32'd1056, 32'd5377, 32'd7918},
{32'd14583, 32'd6270, 32'd10364, 32'd542},
{-32'd10649, 32'd5682, 32'd815, 32'd7353},
{32'd1344, -32'd1894, 32'd2735, -32'd7031},
{32'd5860, 32'd2469, 32'd990, -32'd5504},
{-32'd10199, -32'd2573, -32'd4949, 32'd1159},
{-32'd9926, -32'd799, 32'd2197, 32'd8438},
{-32'd60, -32'd12649, 32'd9016, 32'd6971},
{-32'd6505, -32'd8611, -32'd10821, -32'd4747},
{32'd11978, 32'd4733, -32'd1098, -32'd11259},
{-32'd10048, -32'd2482, 32'd306, -32'd6295},
{32'd4605, -32'd3253, -32'd7567, 32'd14010},
{32'd4112, 32'd3050, 32'd5809, 32'd10525},
{-32'd3152, -32'd11607, -32'd456, -32'd512},
{-32'd6848, 32'd4126, -32'd6535, 32'd8625},
{-32'd1753, 32'd13453, 32'd15887, -32'd6010},
{-32'd9961, -32'd3707, -32'd9860, 32'd7044},
{-32'd8998, -32'd738, -32'd5802, 32'd1283},
{32'd8892, 32'd2981, 32'd3238, 32'd12609},
{32'd4172, 32'd8996, 32'd8821, -32'd8759},
{32'd6596, -32'd194, 32'd8821, -32'd2608},
{32'd3120, -32'd11743, -32'd13772, -32'd552},
{32'd1161, -32'd18046, 32'd2742, -32'd6107},
{-32'd14901, 32'd3465, 32'd134, 32'd1848},
{32'd2210, 32'd8896, -32'd1739, -32'd3158},
{32'd1369, -32'd2875, 32'd1037, -32'd3188},
{32'd500, -32'd16772, 32'd9854, 32'd7600},
{-32'd7839, -32'd8755, -32'd5436, 32'd1406},
{-32'd4883, -32'd355, -32'd3150, -32'd1932},
{-32'd9406, -32'd7827, -32'd1830, 32'd5836},
{-32'd3135, -32'd3958, -32'd1521, 32'd3294},
{-32'd8528, 32'd4529, -32'd1937, -32'd2553},
{-32'd6082, 32'd5130, 32'd6028, -32'd62},
{-32'd5567, -32'd4085, 32'd2355, 32'd3106},
{32'd1261, 32'd207, 32'd1320, 32'd633},
{-32'd6040, 32'd2421, -32'd11888, 32'd18502},
{32'd10107, 32'd10874, -32'd491, 32'd2586},
{-32'd15542, 32'd3613, -32'd894, -32'd13727},
{32'd3306, 32'd8419, -32'd355, 32'd1601},
{-32'd17430, -32'd14515, -32'd4788, 32'd4498},
{32'd10882, -32'd4303, -32'd1628, 32'd2461},
{32'd6579, 32'd936, 32'd1336, -32'd3184},
{32'd236, -32'd14015, -32'd1745, 32'd3374},
{-32'd8342, 32'd3266, 32'd2195, -32'd1785},
{32'd10022, -32'd11304, 32'd262, -32'd5950},
{32'd1800, -32'd190, 32'd5550, -32'd2080},
{32'd853, -32'd1161, -32'd1729, -32'd2093},
{-32'd641, -32'd3493, -32'd3914, -32'd1553},
{-32'd13126, -32'd6137, -32'd3623, -32'd200},
{32'd3962, -32'd2711, -32'd1406, 32'd3841},
{32'd7075, 32'd4073, 32'd2386, 32'd7450},
{32'd15648, -32'd2358, -32'd1832, -32'd6313},
{-32'd6562, -32'd180, -32'd3338, -32'd7373},
{-32'd11555, -32'd8473, 32'd647, -32'd6526},
{-32'd762, 32'd2163, 32'd1853, 32'd7503},
{32'd674, 32'd5801, -32'd14202, 32'd8796},
{-32'd9394, 32'd1053, 32'd3909, -32'd19807},
{-32'd4154, -32'd11729, 32'd3516, 32'd3833},
{32'd16745, 32'd378, 32'd1495, -32'd1019},
{32'd5450, 32'd10578, -32'd9341, -32'd5823},
{-32'd11916, -32'd3025, 32'd4802, 32'd10337},
{32'd11048, -32'd12170, 32'd701, -32'd536},
{32'd17274, -32'd5093, -32'd10171, -32'd2284},
{-32'd11344, 32'd687, -32'd18084, 32'd3825},
{32'd4457, 32'd16225, -32'd14078, -32'd2787},
{-32'd6695, -32'd8475, -32'd10217, 32'd9727},
{32'd11660, -32'd14950, 32'd5726, -32'd10693},
{32'd433, -32'd9182, -32'd1011, 32'd13515},
{-32'd5759, -32'd711, 32'd4699, 32'd8396},
{-32'd1012, -32'd6390, -32'd19058, -32'd256},
{32'd7568, 32'd14136, 32'd9114, 32'd106},
{-32'd2108, -32'd16864, -32'd4014, 32'd21950},
{-32'd7657, -32'd5425, 32'd16112, 32'd2382},
{32'd6344, 32'd3669, 32'd2326, -32'd3083},
{-32'd5760, 32'd333, 32'd8773, 32'd9769},
{32'd6759, 32'd7513, 32'd4338, -32'd3899},
{-32'd1283, -32'd7079, -32'd8844, -32'd905},
{32'd5836, -32'd698, 32'd2518, -32'd4128},
{32'd4634, -32'd5167, -32'd3883, -32'd14274},
{-32'd11965, 32'd5601, 32'd1612, 32'd9384},
{-32'd8359, -32'd4266, 32'd1571, -32'd9704},
{-32'd2422, -32'd5737, 32'd6308, -32'd6811},
{32'd2725, 32'd9947, 32'd596, 32'd5902},
{-32'd2858, -32'd520, 32'd6830, 32'd9340},
{-32'd9532, 32'd3973, 32'd832, 32'd7930},
{-32'd9399, -32'd9750, -32'd10044, 32'd2353},
{-32'd5413, -32'd19690, 32'd16290, 32'd3958},
{32'd3357, 32'd2764, 32'd11054, 32'd4788},
{32'd5471, -32'd4647, 32'd513, 32'd9322},
{-32'd1637, 32'd1653, 32'd10765, -32'd12143},
{-32'd4017, -32'd2076, 32'd8322, 32'd1437},
{32'd1095, 32'd3099, -32'd6201, -32'd2384},
{32'd3752, -32'd3465, 32'd4920, -32'd3191},
{-32'd5895, -32'd1336, 32'd2696, -32'd11750},
{-32'd4330, 32'd3978, -32'd5533, 32'd8206},
{-32'd1132, 32'd7287, 32'd12774, -32'd4124},
{-32'd12502, -32'd6483, 32'd8851, 32'd2230},
{-32'd2570, 32'd22415, 32'd13463, -32'd6492},
{32'd1289, -32'd78, -32'd3242, 32'd3664},
{-32'd4884, -32'd5064, 32'd492, -32'd2720},
{32'd15685, 32'd11478, 32'd4805, -32'd3644},
{-32'd7666, -32'd7837, -32'd12417, -32'd4147},
{-32'd42, -32'd7988, -32'd9572, 32'd14166},
{32'd15566, -32'd13704, 32'd4241, 32'd3096},
{32'd12120, 32'd2886, 32'd3306, 32'd5831},
{32'd12196, 32'd994, 32'd3494, -32'd7487},
{-32'd13105, -32'd16101, -32'd10947, 32'd917},
{32'd3027, 32'd1720, 32'd14599, 32'd1994},
{32'd4848, 32'd7954, -32'd10572, 32'd10851},
{32'd3275, 32'd6232, -32'd10281, 32'd16153},
{32'd9647, 32'd12990, 32'd10924, -32'd5926},
{32'd5042, 32'd8151, -32'd1643, 32'd3265},
{32'd2681, 32'd3519, -32'd1443, 32'd130},
{32'd6466, 32'd5789, 32'd1381, -32'd3497},
{-32'd3403, -32'd4135, 32'd4906, 32'd4864},
{-32'd2919, -32'd11776, -32'd3177, -32'd7411},
{-32'd12282, -32'd2, 32'd2836, -32'd2514},
{-32'd4632, 32'd3731, -32'd11155, -32'd10001},
{32'd10942, -32'd12915, -32'd8750, 32'd1573},
{32'd10610, -32'd2065, -32'd3162, -32'd17522},
{32'd15018, 32'd2947, -32'd4428, -32'd1704},
{-32'd7769, 32'd4991, -32'd1824, 32'd8632},
{-32'd2635, -32'd1268, 32'd219, 32'd1598},
{-32'd269, 32'd10384, 32'd3802, 32'd2997},
{32'd2142, -32'd125, 32'd7125, -32'd783},
{-32'd1206, -32'd1670, -32'd1194, 32'd11662},
{-32'd7913, 32'd6751, 32'd509, 32'd8970},
{-32'd14645, 32'd2676, 32'd5169, 32'd2118},
{32'd7352, 32'd3709, 32'd3731, -32'd2353},
{32'd1326, -32'd4098, -32'd7689, 32'd5557},
{-32'd1038, 32'd7835, 32'd8756, -32'd5701},
{32'd5708, 32'd5692, -32'd4305, -32'd1029},
{-32'd7212, -32'd7527, 32'd3105, -32'd7732},
{32'd8114, -32'd1985, -32'd13263, -32'd5077},
{32'd634, -32'd2344, 32'd4083, -32'd6508},
{-32'd655, -32'd1025, -32'd9417, 32'd7104},
{-32'd1308, 32'd9970, -32'd7325, -32'd7210},
{32'd967, 32'd444, 32'd2020, 32'd6273},
{-32'd15979, 32'd3319, 32'd18309, -32'd369},
{32'd4460, -32'd9331, 32'd12452, 32'd1850},
{-32'd7708, 32'd2250, 32'd6573, 32'd4348},
{-32'd10711, -32'd6714, 32'd9172, 32'd8926},
{32'd7970, -32'd10483, -32'd11252, 32'd11951},
{-32'd4529, 32'd5675, -32'd6164, 32'd5318},
{32'd1496, -32'd1056, -32'd18808, 32'd7898},
{-32'd522, 32'd1152, -32'd1255, -32'd819},
{32'd5172, -32'd3573, -32'd535, -32'd6166},
{-32'd10845, -32'd426, -32'd11471, -32'd5208}
},
{{-32'd12350, 32'd5489, -32'd2955, 32'd8344},
{32'd10249, -32'd6455, -32'd8967, -32'd1763},
{-32'd1684, -32'd1306, 32'd3268, 32'd5385},
{32'd20404, 32'd3114, -32'd5080, -32'd5719},
{32'd10618, 32'd971, -32'd415, -32'd3271},
{-32'd2593, -32'd5126, -32'd3133, 32'd838},
{32'd3422, 32'd2151, 32'd3975, 32'd5966},
{32'd1483, -32'd7135, -32'd3441, -32'd2498},
{32'd12148, -32'd3489, -32'd5632, -32'd1296},
{32'd10114, 32'd6942, 32'd5549, 32'd11190},
{32'd1593, 32'd8062, -32'd9782, -32'd8700},
{-32'd8650, 32'd2286, -32'd1657, -32'd333},
{-32'd4484, -32'd1083, 32'd8626, -32'd6976},
{32'd2256, 32'd5022, -32'd2454, 32'd2774},
{-32'd2741, -32'd6293, -32'd9559, -32'd8029},
{32'd470, 32'd3480, -32'd6728, -32'd1145},
{-32'd716, 32'd2819, 32'd1592, -32'd4045},
{32'd1845, 32'd3646, -32'd6462, 32'd10682},
{32'd10099, 32'd9991, -32'd4439, 32'd6130},
{32'd4949, 32'd10173, -32'd10429, 32'd4349},
{-32'd1014, 32'd5290, -32'd8849, 32'd1655},
{-32'd6964, 32'd11010, 32'd2187, 32'd5349},
{32'd662, 32'd5309, -32'd4230, -32'd4682},
{-32'd11076, 32'd8690, -32'd3448, -32'd642},
{-32'd3529, 32'd11559, 32'd1705, 32'd5084},
{32'd2628, -32'd1829, 32'd724, -32'd2966},
{-32'd6079, -32'd5630, -32'd2102, 32'd5211},
{32'd2513, 32'd8017, 32'd12036, 32'd3956},
{32'd4405, -32'd4479, 32'd9052, 32'd4905},
{-32'd12173, -32'd7690, -32'd7155, -32'd7073},
{-32'd8224, -32'd6854, 32'd8683, -32'd6330},
{32'd6177, -32'd1955, 32'd500, -32'd1955},
{32'd12053, 32'd313, -32'd1416, -32'd4162},
{-32'd815, 32'd657, 32'd1166, -32'd187},
{32'd107, 32'd708, 32'd5726, 32'd5128},
{-32'd8376, 32'd6592, -32'd4755, -32'd3732},
{-32'd3932, -32'd294, -32'd3098, 32'd1017},
{32'd7522, 32'd557, -32'd6701, 32'd2624},
{32'd536, 32'd4460, 32'd729, -32'd2293},
{-32'd6042, -32'd2482, 32'd966, 32'd2005},
{32'd1066, -32'd3453, -32'd5302, 32'd931},
{32'd1090, 32'd13667, 32'd2001, 32'd2955},
{-32'd2277, 32'd9718, 32'd1163, -32'd10918},
{-32'd3051, 32'd4237, 32'd2197, -32'd1121},
{-32'd12985, -32'd8591, -32'd695, 32'd221},
{-32'd3401, -32'd8914, -32'd4951, -32'd6701},
{-32'd10226, -32'd11618, -32'd4053, 32'd7753},
{-32'd19121, -32'd3483, -32'd1978, -32'd261},
{-32'd3853, 32'd8715, -32'd6508, 32'd1450},
{-32'd5126, -32'd2061, -32'd5206, 32'd3214},
{32'd4139, -32'd4063, -32'd2816, -32'd4583},
{32'd1261, 32'd2471, -32'd1563, -32'd1126},
{-32'd1364, 32'd9146, -32'd3765, 32'd1798},
{32'd1241, 32'd1626, 32'd105, -32'd1459},
{-32'd5429, 32'd13141, 32'd2665, 32'd3808},
{32'd3232, -32'd2908, -32'd8164, -32'd2212},
{32'd3146, 32'd1000, -32'd3297, -32'd1398},
{-32'd13519, -32'd743, -32'd1622, -32'd6013},
{32'd3143, -32'd11204, -32'd3937, -32'd4876},
{-32'd11727, -32'd8755, 32'd240, -32'd10861},
{32'd3118, -32'd2110, -32'd1830, -32'd665},
{32'd5577, -32'd236, -32'd525, 32'd2586},
{32'd1393, -32'd168, -32'd4091, -32'd6170},
{32'd621, -32'd4135, -32'd6257, -32'd9087},
{-32'd4786, 32'd12043, -32'd5441, -32'd2799},
{-32'd1105, 32'd7479, 32'd249, 32'd6733},
{32'd480, -32'd5629, 32'd686, 32'd2392},
{-32'd4176, -32'd4142, -32'd4322, 32'd4123},
{-32'd6278, -32'd12203, -32'd12292, 32'd208},
{-32'd2114, -32'd1487, 32'd6616, 32'd2398},
{-32'd4837, 32'd5239, -32'd14510, 32'd5962},
{32'd12737, 32'd3933, 32'd873, 32'd7435},
{-32'd601, -32'd7043, -32'd8084, 32'd6007},
{-32'd8480, -32'd5378, -32'd8463, 32'd6834},
{32'd525, -32'd7664, 32'd5500, 32'd3021},
{-32'd10252, -32'd5522, -32'd4401, -32'd8015},
{-32'd2175, -32'd7152, 32'd1546, 32'd147},
{-32'd9754, -32'd8013, -32'd2756, 32'd2884},
{32'd2287, 32'd5173, 32'd5972, -32'd4010},
{32'd11832, -32'd1319, 32'd6358, -32'd8279},
{32'd3009, -32'd3978, 32'd7871, 32'd3055},
{32'd4660, 32'd10610, 32'd1668, 32'd2226},
{32'd9758, -32'd15129, 32'd1072, -32'd9436},
{32'd6600, -32'd1204, -32'd1805, -32'd5896},
{-32'd3913, -32'd841, 32'd6301, 32'd981},
{-32'd163, 32'd5088, 32'd3149, 32'd5604},
{32'd4805, 32'd11424, -32'd4010, 32'd637},
{-32'd6410, -32'd2430, -32'd6571, -32'd1935},
{32'd846, -32'd10471, 32'd185, -32'd12985},
{-32'd15511, -32'd6396, -32'd1309, -32'd456},
{32'd5489, 32'd3157, 32'd3535, 32'd7083},
{-32'd1934, 32'd8604, -32'd6119, -32'd7375},
{32'd6400, 32'd712, 32'd474, 32'd7820},
{32'd13178, 32'd4578, -32'd5448, 32'd2191},
{32'd7337, 32'd504, 32'd3284, 32'd6104},
{32'd7710, -32'd2400, -32'd5721, -32'd7807},
{-32'd885, 32'd377, 32'd10338, 32'd4356},
{-32'd6086, 32'd1511, 32'd2730, 32'd12515},
{-32'd4759, -32'd5620, 32'd2478, 32'd648},
{32'd6756, -32'd21, 32'd9837, 32'd9299},
{-32'd8255, 32'd11482, -32'd2975, 32'd2372},
{-32'd3201, -32'd5634, 32'd952, 32'd4623},
{-32'd566, -32'd4290, 32'd5134, 32'd7057},
{-32'd2424, -32'd4826, 32'd4069, -32'd4603},
{-32'd986, -32'd4316, -32'd2178, 32'd382},
{-32'd5918, 32'd579, -32'd9512, 32'd1276},
{-32'd7403, -32'd5186, 32'd1204, 32'd7328},
{32'd628, 32'd229, -32'd5678, 32'd42},
{32'd838, 32'd113, 32'd8666, 32'd5183},
{-32'd9728, -32'd8681, -32'd2871, -32'd11833},
{-32'd5920, -32'd5028, -32'd4569, -32'd7599},
{32'd5527, 32'd2054, 32'd1933, -32'd91},
{-32'd2959, 32'd7919, 32'd6365, -32'd7142},
{-32'd585, 32'd12404, -32'd1202, 32'd9499},
{32'd11875, -32'd9910, -32'd926, -32'd698},
{-32'd5746, 32'd1136, -32'd2186, -32'd3715},
{32'd4323, 32'd5598, 32'd11653, -32'd8358},
{32'd1217, 32'd6877, 32'd1849, 32'd8053},
{32'd4731, 32'd7144, -32'd877, -32'd2468},
{32'd8844, 32'd7565, 32'd327, 32'd11024},
{-32'd7401, 32'd9193, 32'd4815, 32'd1030},
{32'd840, 32'd11007, 32'd4516, 32'd4109},
{-32'd11971, -32'd2378, 32'd334, 32'd1917},
{32'd8428, -32'd9373, 32'd1791, -32'd5228},
{32'd8467, 32'd3554, 32'd4616, -32'd8546},
{32'd219, -32'd5841, -32'd421, 32'd555},
{32'd4229, 32'd138, -32'd2851, -32'd8552},
{32'd741, 32'd7848, -32'd5578, -32'd7185},
{32'd4917, -32'd5847, 32'd3616, -32'd10411},
{-32'd5562, -32'd4640, 32'd11692, 32'd2140},
{32'd3039, 32'd1556, -32'd1890, -32'd6736},
{32'd3572, -32'd8968, 32'd813, 32'd3273},
{-32'd10371, -32'd5106, -32'd6669, 32'd1295},
{32'd866, 32'd69, 32'd4821, 32'd4494},
{32'd4298, -32'd1112, 32'd1724, -32'd222},
{32'd192, 32'd1513, -32'd5021, -32'd7855},
{-32'd2441, 32'd1730, -32'd4959, 32'd486},
{-32'd4106, -32'd2476, 32'd3926, -32'd3523},
{32'd16161, 32'd7407, 32'd13067, 32'd5005},
{-32'd3702, -32'd8114, -32'd6068, 32'd2837},
{-32'd3235, 32'd8518, -32'd7540, 32'd11440},
{32'd612, -32'd3189, -32'd1199, -32'd4046},
{-32'd1389, 32'd1728, -32'd6239, -32'd7029},
{32'd9301, 32'd2933, 32'd4439, -32'd9013},
{-32'd3074, 32'd14562, 32'd5735, -32'd359},
{32'd1474, 32'd7358, 32'd760, 32'd2738},
{-32'd10, 32'd6009, -32'd8380, -32'd10103},
{-32'd2200, 32'd7278, 32'd3420, -32'd7895},
{32'd4763, -32'd5051, 32'd4167, 32'd2514},
{-32'd7871, -32'd2983, 32'd4579, 32'd3206},
{-32'd9807, -32'd291, 32'd3123, -32'd6367},
{32'd7215, 32'd4471, -32'd4586, -32'd238},
{-32'd5998, -32'd8398, 32'd419, 32'd794},
{32'd5402, -32'd7677, 32'd6502, -32'd1721},
{-32'd14570, -32'd11300, -32'd5162, -32'd3670},
{32'd7890, -32'd5959, -32'd2769, -32'd7323},
{32'd8119, -32'd3372, 32'd4963, 32'd2981},
{32'd2405, -32'd3573, 32'd3373, -32'd5617},
{-32'd1843, 32'd3279, -32'd830, -32'd5647},
{-32'd8103, 32'd2942, 32'd938, -32'd1524},
{-32'd7310, -32'd1954, -32'd5008, 32'd6069},
{-32'd2652, 32'd6228, 32'd2841, -32'd1390},
{32'd164, -32'd869, -32'd4333, 32'd2054},
{-32'd1803, 32'd4266, 32'd6236, 32'd6037},
{-32'd4820, -32'd3343, 32'd6709, 32'd4621},
{-32'd1767, -32'd1011, -32'd8124, -32'd9458},
{32'd6515, 32'd5526, 32'd3275, 32'd7407},
{32'd2438, 32'd2812, -32'd4977, -32'd7787},
{-32'd6620, -32'd2693, -32'd1474, -32'd10091},
{-32'd11188, 32'd7306, -32'd901, -32'd772},
{-32'd1700, -32'd1211, 32'd4018, 32'd4140},
{32'd9275, -32'd7017, 32'd643, 32'd3181},
{-32'd1076, -32'd1405, 32'd2352, 32'd699},
{32'd1409, 32'd1917, -32'd8059, 32'd6478},
{32'd5252, 32'd1616, 32'd3419, -32'd1024},
{-32'd689, 32'd536, -32'd9626, 32'd1751},
{32'd7810, -32'd1251, 32'd5081, 32'd414},
{32'd1567, -32'd8894, -32'd3182, -32'd8331},
{32'd4911, -32'd955, 32'd1668, 32'd7248},
{32'd3194, -32'd1514, 32'd224, -32'd8886},
{-32'd5779, 32'd5539, -32'd9875, -32'd766},
{32'd4817, -32'd4425, -32'd6735, -32'd1519},
{32'd3693, -32'd98, -32'd15626, -32'd6497},
{-32'd12234, -32'd13746, -32'd1921, -32'd1148},
{-32'd6666, 32'd3520, -32'd315, -32'd397},
{32'd11713, -32'd3509, -32'd9955, -32'd6364},
{32'd5933, -32'd2612, 32'd4968, 32'd2000},
{32'd2547, -32'd1786, -32'd2889, -32'd1561},
{32'd2230, -32'd5541, -32'd3451, -32'd3628},
{-32'd971, -32'd749, 32'd8461, -32'd5307},
{-32'd2191, 32'd3289, -32'd3337, -32'd3042},
{-32'd2407, -32'd2119, -32'd11013, -32'd847},
{-32'd4668, -32'd3629, -32'd10348, -32'd7009},
{32'd8566, 32'd3272, 32'd3282, 32'd6789},
{-32'd4829, -32'd2121, -32'd9174, 32'd10231},
{-32'd5543, 32'd6520, -32'd2544, 32'd3618},
{32'd221, 32'd1751, 32'd1831, 32'd3151},
{-32'd4327, -32'd2437, -32'd7157, -32'd3322},
{32'd3837, -32'd11276, 32'd7111, -32'd7872},
{32'd391, -32'd1138, -32'd1207, 32'd6201},
{-32'd6710, -32'd6014, -32'd6446, -32'd1205},
{32'd11178, -32'd3048, 32'd901, -32'd2260},
{32'd10099, -32'd6575, 32'd5714, 32'd598},
{32'd12932, 32'd738, 32'd521, 32'd10432},
{-32'd15614, -32'd9244, -32'd12548, -32'd866},
{32'd17574, -32'd240, 32'd10037, 32'd2387},
{-32'd3655, 32'd6533, -32'd2717, 32'd2747},
{32'd5115, -32'd7944, 32'd1720, -32'd1776},
{32'd8664, 32'd4551, 32'd5046, -32'd5592},
{32'd5558, -32'd2087, 32'd1332, 32'd4790},
{32'd2583, 32'd2250, 32'd2412, 32'd4266},
{-32'd8283, 32'd9749, -32'd16391, -32'd6721},
{-32'd2963, 32'd10800, 32'd9890, 32'd256},
{32'd1144, -32'd7016, -32'd1602, -32'd70},
{-32'd13360, -32'd7998, -32'd13568, 32'd2909},
{-32'd419, -32'd295, -32'd2289, -32'd6086},
{32'd557, -32'd8276, -32'd6461, 32'd3859},
{-32'd5994, 32'd3969, -32'd4366, -32'd3164},
{32'd10540, 32'd3080, 32'd9607, 32'd798},
{-32'd4106, -32'd7497, 32'd897, 32'd6259},
{-32'd6903, -32'd2251, -32'd10450, -32'd3144},
{32'd2471, 32'd2601, -32'd533, -32'd5043},
{32'd706, -32'd228, 32'd6041, 32'd1273},
{-32'd13983, -32'd1520, 32'd6155, -32'd816},
{-32'd1293, -32'd7918, -32'd3153, 32'd4333},
{32'd4225, -32'd4858, 32'd1761, 32'd3384},
{32'd900, -32'd11252, -32'd4753, -32'd2021},
{-32'd6269, 32'd690, 32'd3806, -32'd2735},
{32'd4118, -32'd2555, 32'd660, -32'd10801},
{32'd2685, 32'd5030, 32'd732, 32'd6980},
{-32'd6296, 32'd3001, -32'd3694, 32'd7797},
{32'd11508, 32'd6333, 32'd3885, -32'd6150},
{32'd1797, 32'd4583, 32'd4461, 32'd1433},
{-32'd1464, -32'd5091, 32'd913, 32'd3913},
{32'd6058, -32'd7329, -32'd451, -32'd1699},
{-32'd605, 32'd540, -32'd7111, -32'd1997},
{32'd1531, -32'd2461, 32'd987, 32'd5161},
{32'd9801, -32'd3402, 32'd6195, -32'd7951},
{-32'd1699, -32'd2394, 32'd6994, -32'd5922},
{32'd31, -32'd1470, -32'd2958, 32'd315},
{-32'd6962, 32'd3497, -32'd8022, 32'd495},
{32'd805, 32'd1, -32'd8890, -32'd3858},
{32'd3045, -32'd7094, -32'd3357, -32'd11057},
{-32'd1231, -32'd9605, -32'd2963, -32'd7545},
{32'd9213, 32'd5878, 32'd3940, 32'd3040},
{-32'd9262, 32'd382, 32'd10399, -32'd3308},
{32'd2854, -32'd14929, 32'd7232, -32'd2462},
{-32'd6971, -32'd1866, -32'd3842, 32'd1382},
{32'd13589, -32'd2308, -32'd8262, 32'd8370},
{32'd3967, -32'd10931, -32'd6312, -32'd11831},
{-32'd132, -32'd494, -32'd13392, -32'd2151},
{32'd675, 32'd2794, 32'd4909, -32'd2155},
{-32'd1697, 32'd6179, 32'd6036, 32'd5325},
{32'd699, 32'd3286, -32'd10415, 32'd3277},
{32'd959, 32'd4928, -32'd9513, 32'd1845},
{32'd4023, 32'd4232, 32'd446, -32'd244},
{32'd5697, 32'd3543, -32'd9388, -32'd5729},
{32'd348, -32'd5543, 32'd5846, 32'd12400},
{-32'd4587, 32'd5363, -32'd3070, -32'd538},
{-32'd732, -32'd4908, 32'd3966, 32'd8326},
{32'd9234, 32'd6571, 32'd6972, 32'd9496},
{-32'd397, 32'd6348, -32'd2506, -32'd1609},
{-32'd6103, -32'd4594, -32'd2474, 32'd2882},
{-32'd7929, -32'd14473, -32'd4849, -32'd1058},
{32'd1288, 32'd2697, 32'd2385, 32'd7485},
{-32'd3163, 32'd2839, 32'd4307, -32'd9150},
{32'd7019, 32'd444, 32'd4159, -32'd7435},
{-32'd1745, 32'd14047, 32'd657, 32'd1693},
{32'd623, -32'd6369, -32'd6257, -32'd10679},
{32'd7404, -32'd756, -32'd384, -32'd10695},
{-32'd6273, -32'd9055, 32'd907, -32'd3213},
{-32'd312, -32'd8586, -32'd3128, 32'd3128},
{-32'd5846, 32'd3794, -32'd4602, 32'd1804},
{-32'd11538, -32'd5468, -32'd159, -32'd4718},
{32'd3683, 32'd6271, -32'd6138, 32'd2692},
{-32'd7695, -32'd441, -32'd4137, -32'd6663},
{32'd6874, 32'd8410, 32'd6748, 32'd7869},
{-32'd3198, -32'd4117, 32'd548, -32'd499},
{-32'd8537, -32'd2544, 32'd10109, -32'd5016},
{32'd1353, -32'd5849, -32'd12515, -32'd71},
{32'd6001, 32'd1852, 32'd6996, 32'd7976},
{32'd6541, 32'd5269, -32'd6298, -32'd14538},
{32'd3240, -32'd1878, -32'd4295, 32'd3679},
{32'd14018, -32'd402, -32'd10888, -32'd75},
{-32'd3933, -32'd1693, 32'd979, -32'd1492},
{-32'd4193, -32'd7975, -32'd6742, -32'd4664},
{32'd1867, -32'd1480, 32'd3971, 32'd1490},
{-32'd6054, 32'd3929, -32'd12336, 32'd3972},
{-32'd8403, 32'd12092, 32'd2258, 32'd2072},
{32'd2250, 32'd3676, 32'd4784, 32'd5290},
{32'd2156, 32'd8753, 32'd4779, -32'd1631},
{32'd5330, 32'd8524, -32'd7236, 32'd2631},
{-32'd861, -32'd6480, -32'd5017, -32'd2883},
{-32'd5317, 32'd491, 32'd4273, 32'd5679},
{32'd2288, -32'd1928, -32'd604, -32'd5955},
{-32'd3648, 32'd564, -32'd4290, -32'd5977},
{-32'd7565, 32'd10723, -32'd742, -32'd5294},
{32'd3146, 32'd2888, 32'd2367, 32'd943},
{-32'd28, -32'd2072, -32'd1877, 32'd417},
{-32'd2745, 32'd4865, -32'd12147, -32'd3450}
},
{{32'd5884, 32'd2868, -32'd2366, 32'd2154},
{-32'd6643, -32'd10989, -32'd992, 32'd14},
{-32'd2673, -32'd3777, -32'd6088, -32'd3188},
{32'd3076, -32'd2840, -32'd3452, -32'd6084},
{-32'd971, 32'd12958, -32'd5515, -32'd2759},
{-32'd2595, 32'd7199, 32'd9258, -32'd7711},
{32'd5773, 32'd10381, -32'd8753, 32'd6402},
{-32'd4221, -32'd4616, -32'd7210, 32'd1464},
{-32'd5614, -32'd4229, -32'd5327, 32'd9281},
{32'd7653, 32'd3949, -32'd2725, -32'd150},
{32'd4862, 32'd2307, 32'd10417, -32'd8524},
{32'd9996, -32'd2521, 32'd307, -32'd15067},
{32'd15894, -32'd8659, 32'd7551, -32'd18522},
{-32'd3817, 32'd1833, -32'd17584, 32'd3858},
{-32'd5991, -32'd736, -32'd6505, 32'd8698},
{32'd9251, -32'd2770, -32'd911, -32'd2675},
{32'd10165, 32'd3714, 32'd820, 32'd1428},
{32'd9084, -32'd9001, 32'd7077, -32'd10133},
{-32'd6084, 32'd3349, -32'd15313, 32'd8650},
{-32'd7048, 32'd573, -32'd3585, -32'd1978},
{-32'd14699, 32'd910, -32'd1750, 32'd11427},
{-32'd14023, -32'd6642, -32'd14164, 32'd1563},
{-32'd7852, -32'd1072, -32'd14130, 32'd6911},
{-32'd843, -32'd8994, 32'd4112, 32'd2209},
{32'd6936, 32'd15958, 32'd7166, 32'd9550},
{-32'd1603, -32'd7249, 32'd4315, 32'd2681},
{-32'd9382, -32'd13157, -32'd3571, 32'd13805},
{32'd67, 32'd11388, 32'd6948, 32'd4663},
{32'd9725, -32'd431, 32'd6679, 32'd6323},
{-32'd3153, 32'd7345, -32'd13983, -32'd8506},
{-32'd4408, 32'd6921, -32'd1417, 32'd7828},
{-32'd8307, -32'd5487, -32'd6786, -32'd6044},
{32'd12226, 32'd290, 32'd8709, -32'd956},
{32'd525, -32'd5338, 32'd9382, -32'd3663},
{32'd7565, 32'd2093, -32'd482, -32'd6776},
{32'd159, -32'd2870, 32'd6384, -32'd8169},
{32'd918, -32'd10095, 32'd7363, 32'd6825},
{32'd10622, 32'd1522, -32'd8669, -32'd1761},
{32'd7479, 32'd13006, 32'd4175, 32'd2538},
{32'd7714, 32'd224, 32'd802, 32'd3750},
{32'd9254, 32'd5774, -32'd4438, -32'd3885},
{32'd8158, 32'd226, -32'd4038, -32'd8448},
{32'd425, -32'd951, -32'd4654, 32'd5367},
{32'd7027, -32'd16012, -32'd7509, 32'd4534},
{-32'd7298, -32'd10769, -32'd7601, -32'd12150},
{32'd6284, -32'd2720, 32'd6702, 32'd5668},
{32'd1186, 32'd1297, -32'd9552, -32'd1068},
{32'd7360, -32'd5053, -32'd7478, -32'd17245},
{-32'd4460, 32'd8558, -32'd1641, -32'd7584},
{-32'd10573, 32'd9447, -32'd5056, 32'd3752},
{-32'd4120, -32'd120, -32'd3979, -32'd5857},
{32'd10901, -32'd348, 32'd13520, -32'd10813},
{32'd423, -32'd8084, -32'd17712, -32'd1012},
{-32'd4444, -32'd6929, 32'd7576, -32'd8650},
{32'd8265, -32'd3113, -32'd2116, 32'd7866},
{-32'd5946, 32'd67, 32'd12297, 32'd6150},
{32'd9102, -32'd2087, -32'd1583, -32'd109},
{32'd527, -32'd1848, -32'd11841, -32'd5485},
{-32'd2073, -32'd5921, -32'd6351, -32'd899},
{-32'd6682, 32'd4798, 32'd11565, 32'd6087},
{-32'd11267, -32'd8401, -32'd2886, 32'd1598},
{32'd6091, 32'd719, 32'd15677, 32'd6783},
{-32'd9618, 32'd2572, -32'd7497, -32'd1232},
{-32'd1193, -32'd9502, -32'd2158, 32'd2253},
{32'd6659, -32'd8852, -32'd9714, 32'd7879},
{32'd5842, 32'd10036, 32'd2634, -32'd3517},
{32'd7126, -32'd10088, 32'd106, 32'd10393},
{-32'd6728, -32'd2025, 32'd2138, 32'd1278},
{32'd4323, -32'd3152, 32'd6045, -32'd6633},
{32'd6616, 32'd4387, -32'd6384, 32'd2573},
{-32'd7638, -32'd2239, 32'd10886, 32'd8009},
{32'd2057, -32'd5667, 32'd6515, 32'd151},
{32'd898, -32'd6803, -32'd1017, -32'd1161},
{-32'd4143, 32'd593, -32'd12768, 32'd3345},
{32'd3068, 32'd1966, 32'd1452, 32'd1535},
{-32'd3602, 32'd8857, -32'd5324, -32'd10737},
{32'd3187, -32'd10748, -32'd1835, -32'd3717},
{-32'd4374, 32'd5905, -32'd8239, 32'd1236},
{-32'd2464, -32'd212, 32'd4098, -32'd238},
{32'd4223, -32'd3044, -32'd5443, -32'd6067},
{32'd4123, -32'd4590, 32'd6966, -32'd6064},
{32'd16070, -32'd4420, -32'd2890, 32'd3481},
{32'd3916, -32'd4861, 32'd9973, 32'd5218},
{32'd4734, 32'd8578, 32'd761, -32'd4917},
{-32'd534, 32'd4627, -32'd2722, -32'd9778},
{32'd3733, 32'd11978, -32'd2386, 32'd8833},
{32'd3129, 32'd5470, -32'd3370, -32'd4101},
{32'd2138, -32'd5311, -32'd330, 32'd3742},
{32'd1293, 32'd9745, 32'd7423, -32'd7526},
{-32'd7760, -32'd4751, -32'd13864, -32'd5260},
{32'd5201, 32'd16652, 32'd9717, -32'd7190},
{-32'd7296, 32'd3598, -32'd9938, 32'd1659},
{32'd1021, 32'd9510, -32'd558, -32'd8559},
{32'd3204, -32'd672, 32'd3418, -32'd10424},
{32'd5117, -32'd2595, 32'd9263, -32'd2094},
{-32'd6738, 32'd486, -32'd1726, -32'd11388},
{32'd10174, 32'd6830, 32'd3310, 32'd434},
{32'd9421, -32'd7332, 32'd642, 32'd2569},
{32'd14836, 32'd1348, -32'd2304, 32'd2213},
{32'd11524, 32'd10526, -32'd4461, -32'd8629},
{32'd1135, -32'd17748, -32'd7253, -32'd6927},
{32'd4741, -32'd6944, -32'd600, -32'd6828},
{32'd14569, 32'd1573, 32'd7790, 32'd2675},
{32'd1307, 32'd8613, -32'd1510, 32'd11784},
{-32'd339, 32'd589, -32'd7421, -32'd4600},
{-32'd9231, 32'd3335, 32'd446, 32'd9203},
{-32'd3002, -32'd3136, -32'd3766, 32'd1245},
{-32'd2089, -32'd5363, 32'd3999, 32'd79},
{32'd3469, -32'd13384, -32'd13367, -32'd12865},
{-32'd14234, -32'd6606, -32'd6652, -32'd5859},
{32'd3296, 32'd6320, 32'd2697, -32'd9742},
{32'd9757, -32'd4918, 32'd3905, 32'd7624},
{-32'd1540, 32'd3592, 32'd6394, 32'd3658},
{-32'd6326, 32'd2202, 32'd4878, -32'd851},
{32'd631, -32'd1007, -32'd14320, 32'd3199},
{-32'd11447, -32'd4751, -32'd16305, 32'd15227},
{32'd8823, 32'd18334, 32'd1413, -32'd5623},
{-32'd7963, -32'd4608, -32'd6182, -32'd412},
{32'd8299, 32'd2108, 32'd1103, 32'd22735},
{32'd4477, 32'd8729, -32'd7017, 32'd2226},
{-32'd3127, 32'd1144, -32'd2221, -32'd3832},
{32'd1014, -32'd5237, -32'd4438, -32'd331},
{32'd2187, 32'd690, 32'd2212, 32'd9610},
{-32'd1868, 32'd10793, -32'd3320, -32'd890},
{32'd5671, 32'd2930, -32'd4230, -32'd4661},
{32'd37, 32'd6770, -32'd723, 32'd3203},
{32'd641, 32'd4990, -32'd6333, 32'd6170},
{-32'd2659, -32'd5246, 32'd9799, 32'd5274},
{-32'd3164, -32'd15122, -32'd12466, -32'd11060},
{-32'd14161, 32'd6257, 32'd5592, 32'd8474},
{-32'd5490, 32'd10122, 32'd2023, 32'd3178},
{32'd1586, 32'd14740, 32'd12125, 32'd1931},
{-32'd16830, -32'd3508, 32'd7466, 32'd1576},
{-32'd950, 32'd13069, -32'd10311, -32'd6342},
{-32'd3568, 32'd3720, 32'd8551, 32'd1970},
{32'd10052, -32'd151, 32'd2240, -32'd6003},
{32'd4548, -32'd4384, 32'd12393, 32'd8501},
{-32'd10271, -32'd15924, 32'd8016, -32'd18092},
{32'd7393, 32'd7345, 32'd5717, 32'd5163},
{32'd3929, -32'd9748, 32'd1595, -32'd5128},
{32'd6918, -32'd4796, -32'd9148, -32'd4179},
{32'd9126, 32'd3863, -32'd3591, -32'd2739},
{32'd4344, 32'd3989, -32'd3044, 32'd10485},
{-32'd2187, 32'd2566, 32'd5713, -32'd374},
{-32'd1155, 32'd3762, 32'd7102, -32'd381},
{-32'd785, 32'd8840, -32'd7062, -32'd2341},
{-32'd8093, -32'd8051, -32'd2992, 32'd2274},
{32'd11387, 32'd596, 32'd10332, 32'd7672},
{-32'd912, -32'd5020, -32'd19229, 32'd2801},
{-32'd6513, -32'd11031, -32'd2600, -32'd892},
{32'd1516, -32'd6672, 32'd1872, 32'd1052},
{-32'd1999, 32'd11713, -32'd8147, -32'd509},
{-32'd3511, -32'd14245, 32'd5102, -32'd122},
{32'd6175, 32'd166, -32'd610, -32'd4365},
{-32'd9830, -32'd1518, 32'd2206, -32'd1191},
{-32'd561, -32'd15654, -32'd1448, 32'd770},
{32'd3243, -32'd8967, -32'd1581, 32'd9763},
{32'd11323, 32'd3456, 32'd7089, 32'd1342},
{32'd8147, -32'd8711, -32'd11536, 32'd6653},
{-32'd3827, -32'd13421, 32'd8865, -32'd9119},
{-32'd16648, -32'd3256, -32'd326, -32'd14514},
{32'd21321, 32'd926, 32'd785, -32'd8927},
{32'd631, -32'd2611, -32'd9061, 32'd544},
{32'd3719, 32'd8296, -32'd1405, -32'd3127},
{-32'd1010, 32'd1630, 32'd14801, 32'd7449},
{-32'd12524, -32'd12559, 32'd12129, 32'd1156},
{-32'd3670, -32'd2910, -32'd7405, -32'd15446},
{-32'd3082, -32'd1063, 32'd6145, 32'd2888},
{32'd3411, -32'd1186, 32'd2812, -32'd12486},
{32'd3839, 32'd617, -32'd5696, 32'd1688},
{-32'd12700, -32'd8441, -32'd5693, -32'd404},
{-32'd8853, -32'd1104, -32'd18, 32'd2435},
{32'd10158, 32'd4766, 32'd6031, -32'd1699},
{-32'd3894, 32'd4354, 32'd831, -32'd7077},
{-32'd6686, 32'd11206, 32'd1613, 32'd1355},
{32'd2625, 32'd2426, -32'd359, -32'd15387},
{32'd4553, 32'd9989, 32'd14366, 32'd12376},
{-32'd500, -32'd1648, 32'd5579, 32'd7684},
{32'd6287, -32'd634, -32'd12701, -32'd3334},
{-32'd2177, -32'd2752, -32'd7016, -32'd10650},
{32'd7898, 32'd26, -32'd4301, -32'd8629},
{32'd2360, 32'd2261, 32'd934, 32'd4077},
{-32'd3950, 32'd188, 32'd530, 32'd9617},
{32'd5402, -32'd5445, -32'd1698, -32'd3405},
{-32'd341, 32'd13792, 32'd3538, -32'd17191},
{-32'd4460, 32'd14945, -32'd832, 32'd13481},
{-32'd5432, 32'd12235, 32'd1580, -32'd2001},
{32'd14591, -32'd5227, -32'd7374, 32'd1289},
{32'd2383, 32'd3218, -32'd6703, 32'd419},
{-32'd2029, 32'd7771, 32'd16625, 32'd469},
{32'd2943, -32'd10245, 32'd4370, -32'd11137},
{-32'd3029, 32'd415, -32'd7485, -32'd176},
{-32'd1710, 32'd7784, -32'd2143, 32'd948},
{-32'd1933, -32'd16118, -32'd5967, 32'd3469},
{32'd733, -32'd16970, -32'd5825, -32'd4074},
{-32'd7067, -32'd15688, -32'd3922, 32'd4914},
{-32'd5834, -32'd11707, -32'd1606, 32'd1038},
{-32'd8743, -32'd8517, 32'd12255, 32'd12170},
{32'd8958, -32'd1406, -32'd16065, 32'd9145},
{32'd4263, -32'd636, 32'd12600, -32'd9090},
{-32'd6866, -32'd4341, -32'd797, 32'd1756},
{32'd7725, 32'd5119, -32'd7268, -32'd8125},
{32'd1845, 32'd6099, 32'd7298, 32'd5418},
{32'd12678, 32'd4896, -32'd136, 32'd5130},
{32'd450, -32'd11027, -32'd14339, -32'd9781},
{32'd869, 32'd4587, 32'd9409, -32'd6135},
{32'd3845, 32'd8572, 32'd4675, 32'd6835},
{-32'd5192, -32'd2004, 32'd16749, 32'd4832},
{32'd4871, 32'd5879, 32'd4587, -32'd11045},
{32'd2616, -32'd5547, 32'd11164, -32'd2733},
{-32'd5915, -32'd3597, -32'd1573, -32'd12426},
{-32'd1294, -32'd1888, 32'd3082, -32'd10689},
{-32'd10848, -32'd11736, -32'd6865, 32'd5510},
{32'd8800, 32'd612, 32'd160, -32'd4297},
{-32'd11293, -32'd4254, -32'd13487, 32'd2073},
{-32'd9346, 32'd8088, -32'd4125, -32'd3918},
{-32'd8480, -32'd1011, 32'd8044, 32'd1600},
{-32'd4148, 32'd502, -32'd9181, 32'd4987},
{32'd4704, -32'd1533, 32'd6902, 32'd14642},
{32'd10076, -32'd13583, -32'd15314, -32'd6017},
{-32'd2961, 32'd7148, 32'd2537, -32'd11828},
{-32'd9482, 32'd2751, 32'd2415, -32'd6130},
{-32'd1239, -32'd7313, -32'd7470, 32'd6930},
{32'd12838, -32'd2764, 32'd9222, 32'd405},
{-32'd4990, 32'd2657, 32'd2903, -32'd3054},
{-32'd6117, -32'd7784, 32'd11808, 32'd3858},
{32'd948, -32'd3001, -32'd9146, -32'd4176},
{-32'd9387, -32'd8906, -32'd10672, 32'd6388},
{-32'd3835, 32'd10603, 32'd5729, 32'd1307},
{32'd14918, -32'd4803, 32'd1910, 32'd2503},
{-32'd18981, -32'd10972, -32'd2502, 32'd5675},
{-32'd1527, 32'd818, -32'd12371, -32'd9826},
{-32'd247, 32'd5443, 32'd1837, 32'd8955},
{-32'd11810, -32'd6355, -32'd14847, -32'd17308},
{32'd4998, 32'd253, -32'd1231, -32'd2417},
{-32'd8946, -32'd4540, -32'd6114, -32'd8027},
{32'd6569, -32'd8409, -32'd3260, 32'd1078},
{32'd1006, -32'd733, 32'd3075, 32'd10508},
{32'd11590, 32'd217, 32'd6795, 32'd4737},
{-32'd4810, -32'd2306, -32'd2249, 32'd2630},
{32'd4872, -32'd14340, -32'd9588, 32'd6148},
{-32'd5908, 32'd2472, 32'd5184, -32'd9669},
{-32'd14753, -32'd15370, -32'd9296, -32'd2205},
{32'd2223, -32'd2376, -32'd830, 32'd2788},
{32'd9448, -32'd122, 32'd11304, 32'd4912},
{32'd6664, -32'd2633, -32'd5352, 32'd6809},
{-32'd1410, -32'd7446, -32'd9776, -32'd9801},
{-32'd1154, -32'd336, 32'd5003, -32'd8951},
{32'd3315, -32'd11284, 32'd112, -32'd4350},
{-32'd3575, -32'd10201, 32'd55, 32'd1426},
{-32'd1857, -32'd10357, 32'd9473, 32'd1698},
{-32'd1708, -32'd4809, -32'd13802, -32'd16491},
{32'd6186, 32'd7184, 32'd3540, -32'd2344},
{-32'd933, 32'd6003, -32'd21787, 32'd1644},
{-32'd3430, -32'd2103, -32'd9115, 32'd7537},
{-32'd3869, -32'd28, 32'd8592, 32'd6991},
{-32'd5010, -32'd8557, -32'd4520, 32'd315},
{32'd1285, 32'd16081, -32'd3799, -32'd4224},
{32'd3372, -32'd15386, 32'd2479, -32'd10919},
{32'd6990, -32'd16740, 32'd6882, 32'd2040},
{32'd4605, -32'd4564, 32'd3413, -32'd5980},
{32'd9247, 32'd214, -32'd7794, -32'd14429},
{-32'd2777, -32'd6922, -32'd9431, -32'd3143},
{32'd362, -32'd6440, -32'd546, -32'd14185},
{32'd3537, 32'd7115, 32'd745, -32'd6988},
{-32'd1270, -32'd4880, -32'd11874, -32'd14357},
{32'd5767, 32'd6446, -32'd1610, -32'd513},
{-32'd2450, -32'd9292, 32'd9096, 32'd8259},
{32'd7126, -32'd6254, 32'd698, -32'd6479},
{-32'd1304, -32'd9784, -32'd6857, 32'd3911},
{-32'd909, 32'd5518, -32'd4904, 32'd9602},
{-32'd9298, 32'd11854, 32'd2693, -32'd603},
{-32'd3388, 32'd5130, -32'd1944, -32'd2630},
{-32'd4090, 32'd2910, -32'd7573, -32'd12023},
{32'd9899, 32'd14704, 32'd2832, -32'd6002},
{-32'd15730, -32'd4659, -32'd5424, 32'd10461},
{32'd12205, 32'd2201, 32'd5244, 32'd2614},
{32'd6945, 32'd5410, 32'd6338, -32'd9277},
{-32'd9915, -32'd13076, -32'd10789, -32'd2176},
{32'd7585, -32'd991, 32'd8635, 32'd6364},
{32'd392, -32'd14278, -32'd13891, 32'd8052},
{32'd4334, 32'd10536, -32'd2347, 32'd921},
{32'd8311, 32'd13451, -32'd3049, 32'd13547},
{-32'd10598, 32'd8467, 32'd5962, 32'd8031},
{-32'd2628, 32'd5948, 32'd2909, 32'd2176},
{-32'd4950, -32'd2679, -32'd1509, 32'd2179},
{-32'd2108, -32'd309, -32'd16514, 32'd8713},
{-32'd754, -32'd18951, -32'd3967, -32'd459},
{-32'd3215, 32'd3390, -32'd8811, 32'd2784},
{32'd3145, 32'd1381, -32'd13398, 32'd1822},
{32'd5590, -32'd18270, 32'd16588, -32'd10666},
{32'd5442, 32'd14316, 32'd16187, 32'd5588},
{32'd2350, 32'd1927, -32'd1912, 32'd7523},
{-32'd8648, 32'd6713, 32'd4791, -32'd12434},
{32'd11202, 32'd6561, 32'd9848, 32'd3426},
{-32'd3875, 32'd2949, 32'd3043, -32'd8330},
{32'd2041, -32'd11957, -32'd2781, -32'd11130},
{32'd3672, -32'd12183, -32'd5788, 32'd113},
{32'd488, 32'd5815, 32'd4433, 32'd10701},
{-32'd5557, -32'd1624, -32'd8720, -32'd1392}
},
{{32'd9800, 32'd7638, 32'd2295, 32'd9853},
{-32'd6006, -32'd3169, -32'd10827, 32'd11313},
{32'd1330, 32'd831, 32'd1524, 32'd10955},
{32'd6768, 32'd14240, 32'd4675, 32'd969},
{-32'd8591, -32'd5564, 32'd12243, 32'd1394},
{-32'd325, -32'd101, 32'd138, -32'd1977},
{-32'd6255, -32'd5346, 32'd3220, -32'd2694},
{-32'd5042, -32'd4196, -32'd4260, 32'd8233},
{32'd3387, -32'd6526, 32'd2817, -32'd1463},
{32'd13252, 32'd9425, 32'd8259, -32'd399},
{32'd321, 32'd846, -32'd13240, -32'd4907},
{-32'd8615, 32'd2951, -32'd3666, 32'd3921},
{32'd6814, 32'd4418, 32'd2824, 32'd64},
{-32'd784, -32'd4437, 32'd3266, -32'd6704},
{-32'd6091, -32'd779, 32'd544, -32'd4169},
{32'd569, 32'd4600, 32'd3720, -32'd4248},
{-32'd4974, 32'd5422, -32'd5198, -32'd4344},
{32'd1413, 32'd1250, -32'd5966, 32'd5059},
{32'd2074, -32'd5032, -32'd9322, -32'd6317},
{-32'd6743, 32'd1189, -32'd5287, 32'd2268},
{32'd6021, -32'd3341, 32'd2069, -32'd666},
{-32'd1279, -32'd3373, -32'd10144, 32'd7823},
{-32'd12515, -32'd9003, -32'd564, -32'd1487},
{32'd7810, -32'd15526, -32'd9400, -32'd442},
{32'd10226, 32'd5669, -32'd3041, -32'd3924},
{32'd3030, -32'd4663, -32'd4571, 32'd6626},
{32'd4089, 32'd1586, -32'd2443, 32'd1313},
{32'd4569, 32'd752, -32'd441, -32'd1961},
{32'd4202, 32'd237, -32'd2311, -32'd1929},
{-32'd2088, -32'd9128, -32'd1782, -32'd2273},
{32'd2678, -32'd64, 32'd4956, 32'd5574},
{-32'd8783, -32'd13086, -32'd18285, 32'd2250},
{32'd6283, 32'd7155, 32'd2709, -32'd665},
{32'd4584, -32'd5242, -32'd2856, -32'd1292},
{32'd11298, 32'd6605, 32'd6230, -32'd6281},
{32'd3851, -32'd6660, -32'd6497, 32'd3614},
{-32'd19086, -32'd5187, -32'd1867, -32'd855},
{32'd935, 32'd5263, 32'd12169, -32'd10127},
{-32'd3078, 32'd8231, -32'd5716, 32'd769},
{32'd3001, -32'd2219, -32'd15383, -32'd8093},
{32'd10124, -32'd2672, -32'd1570, 32'd3717},
{32'd5034, -32'd4086, 32'd7428, 32'd4718},
{-32'd1966, -32'd4865, -32'd1037, 32'd8259},
{-32'd428, -32'd2753, -32'd4357, -32'd3857},
{-32'd3113, -32'd10528, -32'd5604, -32'd3493},
{32'd11771, 32'd10009, -32'd2959, -32'd4392},
{-32'd931, 32'd2441, 32'd43, 32'd5682},
{-32'd6305, -32'd1501, -32'd6824, 32'd3393},
{-32'd5487, 32'd7982, 32'd5597, 32'd4255},
{-32'd14089, -32'd4393, 32'd1546, 32'd574},
{-32'd5907, -32'd10133, 32'd5242, 32'd10989},
{32'd341, 32'd7356, 32'd5179, -32'd756},
{32'd7844, -32'd3489, -32'd8545, 32'd7843},
{32'd5271, 32'd2301, -32'd6958, 32'd3140},
{32'd5145, 32'd2315, 32'd7652, -32'd2352},
{-32'd8167, -32'd5043, -32'd4263, 32'd3125},
{-32'd1255, 32'd13759, 32'd5440, -32'd7040},
{32'd1067, -32'd2565, -32'd7844, -32'd3283},
{-32'd2613, -32'd1983, -32'd6020, -32'd4465},
{-32'd952, 32'd2222, 32'd6360, 32'd1026},
{-32'd14200, -32'd6646, 32'd622, 32'd1855},
{-32'd1006, 32'd205, -32'd150, -32'd12928},
{-32'd3559, -32'd9326, -32'd5148, 32'd2356},
{-32'd1132, -32'd6302, -32'd2691, 32'd5527},
{32'd1915, 32'd2167, 32'd627, -32'd726},
{32'd11418, 32'd9336, 32'd2141, 32'd549},
{-32'd1554, 32'd1421, -32'd10852, 32'd540},
{-32'd13768, -32'd15084, 32'd435, -32'd1838},
{32'd5423, 32'd302, 32'd848, 32'd13904},
{32'd1433, -32'd2245, 32'd2805, 32'd13309},
{32'd5340, -32'd4653, 32'd762, 32'd4268},
{32'd975, -32'd5421, -32'd4277, 32'd2548},
{32'd2042, 32'd103, -32'd5768, 32'd11887},
{-32'd6340, -32'd1834, -32'd5485, 32'd714},
{32'd3872, 32'd2605, 32'd7961, 32'd31},
{32'd10401, 32'd4501, 32'd1329, 32'd477},
{32'd555, -32'd533, 32'd6771, -32'd11070},
{-32'd12818, 32'd6614, 32'd300, -32'd3340},
{32'd9546, -32'd2536, 32'd4067, 32'd1958},
{-32'd1951, 32'd1518, 32'd3084, 32'd3174},
{-32'd5228, -32'd174, 32'd17322, -32'd4543},
{32'd11371, 32'd17438, 32'd776, 32'd8626},
{-32'd5855, -32'd5148, -32'd12121, 32'd4799},
{-32'd4366, 32'd8493, -32'd12445, -32'd7693},
{-32'd3555, -32'd6960, -32'd8515, 32'd10150},
{-32'd5485, -32'd8962, -32'd5960, 32'd9551},
{32'd6045, -32'd291, -32'd3372, 32'd6324},
{-32'd6309, -32'd7360, -32'd1454, 32'd661},
{-32'd1629, -32'd1180, 32'd3694, 32'd231},
{-32'd1065, -32'd1396, 32'd4917, 32'd6674},
{32'd6589, 32'd3419, -32'd1874, -32'd8437},
{-32'd5997, -32'd4188, -32'd678, 32'd4677},
{32'd7488, 32'd4693, 32'd10091, 32'd3480},
{-32'd5298, -32'd9272, 32'd4248, -32'd6912},
{-32'd2104, 32'd2516, -32'd7854, 32'd691},
{32'd3240, 32'd2691, -32'd1820, 32'd295},
{32'd1664, -32'd743, 32'd4554, -32'd2381},
{-32'd7600, -32'd14564, 32'd7690, -32'd2697},
{-32'd11509, -32'd2798, -32'd8851, -32'd637},
{32'd10009, 32'd5225, 32'd2850, -32'd2124},
{32'd2529, -32'd4587, -32'd4313, -32'd7460},
{32'd2467, -32'd8023, -32'd1306, 32'd1949},
{32'd2591, -32'd2856, -32'd3344, -32'd6787},
{32'd8084, 32'd10141, 32'd4035, -32'd7497},
{32'd3283, 32'd3326, 32'd4720, -32'd2717},
{-32'd7188, -32'd7765, 32'd7144, 32'd1959},
{-32'd8284, -32'd5578, -32'd4558, 32'd2430},
{32'd3510, 32'd1139, 32'd103, -32'd2223},
{32'd7566, 32'd18325, 32'd5866, -32'd6506},
{-32'd7305, -32'd9154, -32'd323, -32'd2271},
{-32'd6284, -32'd6090, 32'd3276, -32'd5524},
{32'd5471, -32'd481, -32'd2948, -32'd836},
{-32'd7227, 32'd5119, 32'd4458, -32'd4136},
{32'd7484, 32'd3936, 32'd138, -32'd3684},
{-32'd9680, -32'd9755, 32'd1148, 32'd4035},
{-32'd12869, -32'd11682, -32'd4826, 32'd5800},
{-32'd9228, -32'd10060, -32'd5166, 32'd5585},
{-32'd5879, -32'd4614, -32'd1353, -32'd14189},
{32'd9172, 32'd5606, 32'd278, 32'd243},
{32'd4514, 32'd11677, 32'd4555, 32'd2884},
{-32'd11398, 32'd7470, -32'd475, -32'd694},
{32'd7769, 32'd3357, 32'd1049, -32'd4621},
{-32'd6729, 32'd2134, 32'd4836, 32'd6914},
{32'd2097, 32'd8004, -32'd9267, 32'd2450},
{-32'd4433, 32'd10826, -32'd5195, 32'd8625},
{-32'd553, -32'd1929, 32'd682, -32'd9544},
{-32'd5007, -32'd10938, -32'd3043, -32'd495},
{32'd1247, -32'd6058, -32'd11010, -32'd7193},
{32'd698, -32'd14131, -32'd9512, -32'd6978},
{-32'd2640, -32'd2591, 32'd2317, -32'd3074},
{-32'd5809, -32'd3869, 32'd1691, 32'd10681},
{-32'd9233, -32'd9997, -32'd3823, 32'd3101},
{-32'd5440, 32'd2695, -32'd11934, -32'd5316},
{-32'd4301, -32'd5285, 32'd1745, 32'd3469},
{32'd4080, -32'd3263, 32'd6646, 32'd3230},
{-32'd1169, -32'd3138, -32'd4918, 32'd255},
{-32'd403, 32'd13822, 32'd748, 32'd1911},
{32'd3404, 32'd918, -32'd268, 32'd5360},
{32'd10858, 32'd3129, 32'd3639, 32'd1717},
{-32'd13233, -32'd5674, -32'd1576, 32'd9973},
{-32'd7828, -32'd3136, -32'd5301, -32'd926},
{-32'd67, 32'd379, -32'd4218, 32'd3154},
{32'd6878, 32'd1972, -32'd7600, 32'd9786},
{32'd163, -32'd1044, -32'd772, -32'd6081},
{32'd9426, 32'd1088, -32'd1660, -32'd864},
{-32'd5892, -32'd1797, 32'd8512, 32'd10681},
{32'd2129, -32'd4662, 32'd1611, -32'd6369},
{-32'd786, 32'd505, -32'd7066, -32'd8952},
{32'd10274, 32'd80, 32'd3678, 32'd705},
{-32'd14582, -32'd3314, -32'd7766, 32'd9133},
{-32'd10047, -32'd1399, 32'd2422, -32'd5556},
{32'd6360, 32'd12961, 32'd10082, -32'd12955},
{-32'd835, -32'd834, 32'd1900, -32'd4803},
{32'd11577, -32'd598, -32'd6083, -32'd7636},
{-32'd5753, -32'd2314, -32'd5089, -32'd5900},
{-32'd5613, 32'd1851, -32'd823, -32'd1236},
{-32'd2791, 32'd7921, 32'd3623, 32'd3074},
{-32'd8170, 32'd7714, 32'd2946, -32'd9540},
{-32'd2309, -32'd732, -32'd601, 32'd4435},
{32'd0, -32'd4581, 32'd1975, 32'd6785},
{-32'd4483, -32'd2514, -32'd358, 32'd16913},
{-32'd1025, 32'd2914, 32'd12829, -32'd5906},
{-32'd6907, -32'd6927, -32'd2358, -32'd6298},
{32'd10882, 32'd2194, 32'd3849, -32'd2275},
{32'd3149, 32'd3604, 32'd3013, -32'd2909},
{32'd1882, 32'd902, -32'd4158, -32'd1379},
{-32'd13902, 32'd9519, -32'd5031, -32'd4463},
{32'd1826, -32'd4006, -32'd13409, 32'd5831},
{32'd5728, 32'd8329, 32'd882, 32'd1628},
{-32'd7407, 32'd1445, 32'd15385, 32'd1073},
{32'd1572, -32'd1869, -32'd2210, -32'd10473},
{32'd92, 32'd2396, -32'd15177, -32'd1380},
{32'd13366, 32'd11063, -32'd123, -32'd6777},
{-32'd7318, -32'd2947, -32'd160, -32'd12817},
{-32'd206, 32'd1090, 32'd6577, 32'd285},
{32'd9651, 32'd2978, 32'd1033, -32'd7188},
{32'd3281, 32'd2501, 32'd5534, -32'd3948},
{32'd3340, -32'd1943, -32'd2354, 32'd936},
{32'd3643, -32'd1266, 32'd2430, -32'd928},
{-32'd3934, -32'd11151, -32'd7052, -32'd7296},
{-32'd1313, -32'd1109, -32'd4690, 32'd925},
{-32'd3079, 32'd879, -32'd2981, -32'd3405},
{-32'd798, 32'd2477, -32'd5494, -32'd1524},
{32'd8755, -32'd3858, 32'd1791, -32'd523},
{32'd1564, -32'd1142, -32'd5980, -32'd3049},
{32'd1704, 32'd153, 32'd255, -32'd1313},
{32'd10658, 32'd282, -32'd3706, 32'd8605},
{32'd2035, -32'd15006, -32'd4515, -32'd3609},
{32'd5058, -32'd2525, 32'd5565, -32'd6982},
{-32'd1263, 32'd1680, -32'd11777, 32'd8005},
{-32'd1422, -32'd4257, 32'd1225, 32'd4182},
{-32'd5109, 32'd1743, -32'd9000, -32'd6658},
{32'd6100, -32'd3684, -32'd6160, -32'd4880},
{32'd6995, 32'd2406, -32'd1665, 32'd3221},
{-32'd310, -32'd238, 32'd6574, 32'd3613},
{32'd5944, -32'd6111, -32'd1283, 32'd2302},
{32'd11247, -32'd122, 32'd4722, -32'd6353},
{32'd5035, 32'd8309, 32'd6625, 32'd1786},
{32'd5793, -32'd4679, 32'd2440, 32'd11283},
{32'd2125, 32'd3818, 32'd3202, -32'd8006},
{-32'd10849, -32'd8708, -32'd7903, 32'd1288},
{-32'd4486, -32'd10332, -32'd5441, -32'd7920},
{32'd1621, -32'd11807, -32'd2708, -32'd1472},
{-32'd3227, 32'd1809, 32'd1791, 32'd963},
{-32'd14867, -32'd806, -32'd5890, 32'd2143},
{32'd2450, 32'd3700, -32'd10856, -32'd4347},
{32'd3004, -32'd8393, -32'd6451, 32'd2931},
{-32'd9880, -32'd5877, -32'd4809, -32'd6},
{32'd5223, 32'd8744, 32'd10286, 32'd2372},
{32'd3537, 32'd6223, 32'd173, -32'd3818},
{-32'd2991, -32'd5423, -32'd1530, -32'd3031},
{-32'd3646, 32'd1620, 32'd6247, -32'd4957},
{-32'd2642, -32'd6812, -32'd5313, 32'd19781},
{32'd13832, -32'd2314, 32'd5929, -32'd6367},
{-32'd9227, 32'd3509, 32'd6851, -32'd13529},
{-32'd7271, -32'd18885, -32'd10484, -32'd4504},
{32'd4074, -32'd10708, -32'd5015, 32'd1952},
{32'd4214, 32'd4209, 32'd249, 32'd1141},
{-32'd1666, -32'd2648, 32'd7537, -32'd9614},
{-32'd1738, -32'd1041, 32'd4608, 32'd3625},
{-32'd5959, -32'd2027, -32'd10203, -32'd6160},
{32'd1926, -32'd4661, 32'd3525, 32'd5240},
{-32'd6578, 32'd1212, 32'd13700, -32'd5561},
{32'd7777, 32'd3427, 32'd2066, -32'd1953},
{-32'd1168, -32'd2478, 32'd1775, 32'd6247},
{-32'd3206, -32'd5605, 32'd4219, 32'd3642},
{-32'd3507, -32'd4938, -32'd6360, 32'd942},
{-32'd3331, -32'd6843, 32'd2177, -32'd757},
{-32'd7207, -32'd367, 32'd2971, 32'd7856},
{32'd1113, 32'd9033, -32'd11772, 32'd2311},
{-32'd2906, -32'd10261, -32'd4420, 32'd191},
{-32'd6850, 32'd1373, -32'd50, -32'd7804},
{32'd5870, -32'd5946, 32'd8879, 32'd12074},
{-32'd3168, -32'd5032, 32'd7588, 32'd0},
{-32'd5967, 32'd2502, -32'd11646, -32'd2630},
{32'd3938, -32'd8162, -32'd9261, 32'd1013},
{-32'd2736, -32'd49, -32'd2293, -32'd8933},
{32'd11649, 32'd2320, 32'd5510, 32'd2750},
{32'd8910, 32'd6024, 32'd4369, -32'd10587},
{-32'd6877, -32'd3253, 32'd1146, 32'd5531},
{-32'd7711, 32'd5465, -32'd7576, 32'd7112},
{-32'd5865, -32'd4610, 32'd1753, 32'd3497},
{-32'd9148, -32'd2531, 32'd1477, 32'd4642},
{-32'd3615, -32'd340, -32'd2872, -32'd1211},
{32'd8913, 32'd7192, 32'd10014, -32'd2465},
{32'd3344, 32'd5863, 32'd8797, -32'd150},
{32'd5, -32'd1113, -32'd1303, 32'd2815},
{32'd3305, -32'd1853, -32'd6457, 32'd2265},
{32'd11474, -32'd6143, 32'd5217, 32'd5054},
{32'd1642, -32'd1600, 32'd2506, -32'd1839},
{-32'd4189, -32'd9354, -32'd6286, 32'd811},
{32'd2030, 32'd6570, 32'd1367, -32'd3796},
{-32'd939, 32'd3685, 32'd4222, -32'd9583},
{32'd11904, -32'd2473, 32'd5169, -32'd800},
{-32'd3838, -32'd8689, -32'd10648, -32'd9279},
{32'd757, 32'd5850, -32'd4840, 32'd7114},
{-32'd8504, -32'd27, -32'd130, -32'd9743},
{32'd1021, -32'd3272, 32'd3325, 32'd5305},
{-32'd1753, 32'd2661, -32'd6775, -32'd13816},
{-32'd2003, 32'd3370, 32'd3390, -32'd4381},
{32'd3300, -32'd750, -32'd9594, -32'd1377},
{32'd7759, 32'd3404, -32'd285, 32'd5869},
{-32'd2784, -32'd4400, -32'd1174, 32'd2128},
{-32'd13625, 32'd9095, 32'd3800, 32'd289},
{-32'd4170, -32'd4468, 32'd6932, -32'd9120},
{32'd9130, 32'd7361, -32'd4740, 32'd7128},
{-32'd3256, 32'd2949, 32'd901, 32'd2143},
{-32'd4732, -32'd7815, -32'd2809, -32'd663},
{32'd11195, 32'd887, -32'd6804, -32'd271},
{32'd9628, -32'd6332, -32'd1128, -32'd1543},
{-32'd1174, 32'd3166, 32'd8233, -32'd5060},
{32'd504, 32'd13959, -32'd2225, 32'd8603},
{-32'd2336, -32'd8504, -32'd2483, 32'd2714},
{32'd2206, -32'd13031, 32'd1742, 32'd833},
{32'd1415, 32'd4937, -32'd982, -32'd5694},
{-32'd1074, -32'd9205, -32'd6477, -32'd1499},
{32'd13848, 32'd8702, 32'd8703, 32'd1984},
{32'd14590, 32'd4585, 32'd6713, -32'd6643},
{-32'd4238, -32'd5806, 32'd3726, -32'd1629},
{-32'd4962, 32'd26, -32'd11888, 32'd4401},
{32'd10551, 32'd774, -32'd147, 32'd12143},
{32'd8778, 32'd9124, 32'd1077, 32'd10390},
{-32'd9759, -32'd102, 32'd4505, 32'd5173},
{32'd9183, -32'd4514, 32'd543, 32'd7828},
{-32'd2909, 32'd4436, 32'd6941, -32'd1431},
{-32'd719, -32'd1013, -32'd6786, -32'd1122},
{-32'd2275, 32'd1506, 32'd1332, 32'd434},
{-32'd1750, -32'd1612, -32'd5110, -32'd3062},
{-32'd3762, 32'd2645, 32'd10364, 32'd4962},
{-32'd399, 32'd700, -32'd3113, 32'd5113},
{-32'd520, -32'd12600, 32'd7030, 32'd987},
{32'd705, 32'd3121, 32'd3710, -32'd253},
{32'd4117, 32'd4729, 32'd869, 32'd5723},
{32'd3944, -32'd3515, 32'd315, -32'd2167},
{-32'd274, -32'd3153, -32'd569, 32'd1040},
{-32'd9523, -32'd403, -32'd713, -32'd4234},
{-32'd2339, -32'd520, -32'd9823, -32'd5517},
{32'd6844, 32'd12653, 32'd4162, 32'd7346},
{32'd977, 32'd1672, 32'd6946, -32'd78},
{-32'd4748, -32'd2104, -32'd4229, 32'd952}
},
{{-32'd7736, 32'd6630, 32'd4631, 32'd6500},
{-32'd6999, -32'd6335, -32'd2325, -32'd900},
{32'd259, 32'd3579, 32'd4279, -32'd210},
{32'd16697, 32'd9133, 32'd6698, 32'd16027},
{-32'd3025, 32'd3326, -32'd1314, 32'd2283},
{32'd247, 32'd275, 32'd2961, 32'd8851},
{-32'd8810, -32'd779, 32'd8658, 32'd5126},
{-32'd822, -32'd400, 32'd4934, 32'd4377},
{32'd1569, 32'd6896, 32'd3496, -32'd4138},
{32'd4029, 32'd6116, 32'd4413, 32'd7120},
{-32'd7185, 32'd1508, -32'd4334, -32'd5151},
{32'd9436, 32'd3079, 32'd1635, 32'd561},
{32'd5687, -32'd1853, -32'd1309, -32'd1828},
{-32'd3431, -32'd3814, -32'd1031, 32'd4198},
{-32'd6877, 32'd3934, -32'd1836, -32'd1580},
{32'd10738, -32'd142, 32'd965, -32'd6841},
{-32'd8621, 32'd1408, 32'd2583, -32'd4553},
{32'd4970, 32'd4971, -32'd1039, -32'd4329},
{-32'd7249, -32'd1028, -32'd3640, 32'd4620},
{-32'd2123, 32'd5776, -32'd3464, -32'd2682},
{32'd1160, -32'd2313, 32'd752, 32'd107},
{-32'd6881, -32'd3059, -32'd6989, -32'd4589},
{32'd642, 32'd2035, -32'd8769, 32'd1252},
{-32'd4357, -32'd4557, -32'd8943, -32'd5147},
{32'd385, 32'd3098, -32'd2591, 32'd8792},
{32'd12346, 32'd2620, 32'd13649, 32'd7144},
{-32'd8512, 32'd3834, -32'd793, -32'd1158},
{32'd9392, -32'd66, 32'd4983, -32'd7502},
{32'd2247, 32'd6438, -32'd83, -32'd7072},
{-32'd1717, 32'd7041, -32'd9567, -32'd4560},
{-32'd1124, 32'd1468, 32'd4397, -32'd2305},
{-32'd9717, -32'd3835, -32'd5887, -32'd8229},
{-32'd1444, 32'd897, -32'd618, 32'd7602},
{32'd8137, 32'd836, -32'd5157, 32'd2712},
{-32'd1556, 32'd6239, 32'd5536, 32'd4580},
{-32'd7859, 32'd4163, -32'd2692, -32'd8598},
{-32'd7678, -32'd2916, 32'd4988, 32'd4879},
{-32'd9661, 32'd5835, 32'd1522, 32'd3305},
{32'd4826, 32'd373, 32'd4576, -32'd5548},
{-32'd14748, -32'd3190, -32'd6611, -32'd3680},
{-32'd5110, -32'd4168, -32'd6983, -32'd4451},
{-32'd1848, 32'd4890, -32'd2220, -32'd2504},
{-32'd3483, 32'd413, 32'd507, 32'd2663},
{-32'd622, -32'd5065, -32'd4419, 32'd584},
{32'd3462, -32'd1470, -32'd777, -32'd10569},
{32'd5816, -32'd3238, -32'd3283, -32'd1714},
{-32'd5309, -32'd276, -32'd8322, -32'd409},
{-32'd11177, -32'd507, 32'd681, 32'd543},
{32'd560, 32'd9506, 32'd1610, 32'd2637},
{-32'd5777, -32'd524, -32'd1720, 32'd6008},
{-32'd3032, 32'd3714, -32'd1274, -32'd5192},
{-32'd3664, -32'd3111, 32'd3760, 32'd4963},
{-32'd9773, 32'd3344, 32'd334, 32'd5215},
{-32'd5582, 32'd3378, -32'd6157, 32'd3640},
{32'd839, -32'd751, 32'd1083, -32'd3614},
{32'd4607, -32'd2073, 32'd1219, -32'd3314},
{32'd2389, 32'd5936, 32'd12039, 32'd1223},
{32'd3067, 32'd6402, -32'd7524, 32'd772},
{-32'd12141, -32'd2881, -32'd7834, 32'd5879},
{-32'd13266, 32'd4913, 32'd3259, -32'd3078},
{-32'd6519, 32'd332, 32'd2170, 32'd9582},
{-32'd704, -32'd7933, -32'd1021, 32'd8953},
{-32'd11128, 32'd1736, -32'd5847, -32'd5298},
{-32'd535, 32'd8380, 32'd3195, -32'd2366},
{-32'd1836, 32'd624, 32'd807, 32'd1072},
{32'd12899, 32'd7053, 32'd7607, 32'd10536},
{32'd9831, -32'd1334, -32'd1770, -32'd3716},
{32'd4562, 32'd1220, 32'd3593, -32'd6154},
{-32'd8767, 32'd7565, -32'd4661, -32'd3722},
{32'd6860, -32'd1899, 32'd536, -32'd3227},
{-32'd1528, -32'd7140, 32'd2057, -32'd9142},
{32'd3981, -32'd80, -32'd359, -32'd3328},
{-32'd3306, -32'd6024, -32'd6076, -32'd15176},
{32'd1696, 32'd10853, 32'd700, 32'd3487},
{32'd6966, 32'd10761, 32'd8282, -32'd7297},
{32'd5448, -32'd412, 32'd6846, 32'd2721},
{32'd902, -32'd8644, -32'd4577, 32'd7447},
{-32'd4508, 32'd2413, 32'd2396, -32'd291},
{32'd3299, 32'd1222, 32'd5731, 32'd1571},
{32'd9860, -32'd3128, 32'd4387, 32'd2302},
{-32'd10023, 32'd6571, 32'd6030, 32'd1338},
{-32'd2973, 32'd5346, 32'd1595, -32'd4730},
{-32'd2997, -32'd1422, -32'd2322, -32'd10686},
{-32'd8603, -32'd6762, 32'd4962, -32'd6045},
{32'd2583, -32'd4308, -32'd8031, -32'd7636},
{-32'd3670, -32'd3601, -32'd892, -32'd7584},
{-32'd533, 32'd4113, 32'd15076, 32'd7209},
{-32'd9119, -32'd7157, -32'd7492, -32'd8904},
{32'd7227, 32'd6240, -32'd462, 32'd1893},
{-32'd11201, 32'd1202, -32'd124, 32'd761},
{-32'd3676, 32'd4307, 32'd2391, 32'd1400},
{-32'd3030, -32'd20, -32'd8668, -32'd5586},
{32'd5624, 32'd379, 32'd1058, 32'd8294},
{32'd13414, 32'd5185, 32'd5471, 32'd3594},
{32'd10951, 32'd339, 32'd3983, 32'd3819},
{-32'd5087, -32'd1267, -32'd596, -32'd4702},
{32'd1613, 32'd602, 32'd8522, 32'd3441},
{32'd7651, 32'd1752, 32'd7180, 32'd1812},
{-32'd5115, 32'd5049, -32'd3470, -32'd4676},
{32'd3049, 32'd3425, -32'd366, 32'd11202},
{32'd99, -32'd4402, 32'd4648, 32'd4643},
{-32'd11270, 32'd1171, -32'd4471, -32'd8898},
{32'd4246, -32'd8227, 32'd1598, 32'd2661},
{-32'd6630, -32'd4500, 32'd3146, -32'd208},
{32'd12803, -32'd7364, -32'd1236, 32'd471},
{32'd11269, 32'd5682, 32'd919, 32'd1809},
{32'd1038, -32'd3174, 32'd2399, -32'd666},
{32'd10820, -32'd1520, -32'd1853, 32'd3322},
{-32'd2928, 32'd386, 32'd1823, 32'd8901},
{-32'd5991, -32'd4590, 32'd381, 32'd2721},
{-32'd1813, -32'd4992, 32'd4305, 32'd593},
{-32'd3983, 32'd3657, -32'd7093, -32'd4476},
{-32'd317, 32'd892, 32'd374, -32'd7175},
{32'd80, 32'd5063, 32'd7437, 32'd1168},
{32'd4975, 32'd2707, -32'd535, 32'd3671},
{-32'd5331, -32'd2887, 32'd5245, -32'd7587},
{32'd2440, 32'd5834, 32'd7129, -32'd2129},
{-32'd1934, -32'd8244, 32'd1601, -32'd4622},
{-32'd1445, -32'd4147, 32'd5960, -32'd10714},
{-32'd6107, 32'd6721, 32'd2657, 32'd9979},
{-32'd1487, 32'd6751, 32'd633, -32'd737},
{-32'd6718, -32'd4096, -32'd815, 32'd2225},
{32'd12017, 32'd1165, -32'd10136, 32'd2413},
{32'd2077, -32'd199, -32'd2865, -32'd5608},
{32'd5601, 32'd4129, -32'd734, -32'd161},
{-32'd4532, -32'd1498, 32'd5664, 32'd7987},
{-32'd5482, -32'd2080, -32'd2457, 32'd1109},
{-32'd1885, -32'd380, 32'd3872, -32'd2769},
{-32'd9317, -32'd7634, -32'd4079, -32'd26},
{-32'd8407, -32'd5659, 32'd2394, 32'd3590},
{-32'd3264, 32'd2023, 32'd4639, -32'd8042},
{-32'd11989, -32'd16341, -32'd375, -32'd9745},
{-32'd6569, -32'd4080, 32'd6141, 32'd1911},
{32'd4328, 32'd396, -32'd551, 32'd5204},
{32'd8119, -32'd2581, -32'd3323, -32'd9013},
{32'd1457, 32'd3903, -32'd9107, -32'd6134},
{32'd7275, -32'd5261, -32'd4500, -32'd6798},
{32'd8103, -32'd4331, 32'd2565, -32'd3752},
{32'd1364, -32'd75, 32'd1628, -32'd5167},
{-32'd11786, -32'd3450, -32'd3173, 32'd6737},
{-32'd5530, -32'd298, -32'd548, -32'd3011},
{-32'd4610, -32'd2184, 32'd3092, 32'd2419},
{32'd2099, -32'd5761, -32'd6314, -32'd133},
{-32'd5639, 32'd1949, -32'd3551, -32'd2772},
{-32'd7466, -32'd416, 32'd4099, -32'd1448},
{32'd3727, 32'd2843, 32'd8870, 32'd8376},
{32'd185, 32'd8018, -32'd884, -32'd10646},
{-32'd5413, -32'd7303, -32'd5736, -32'd3073},
{32'd1861, 32'd3962, 32'd9655, 32'd7501},
{-32'd1605, 32'd3743, 32'd7349, 32'd4651},
{-32'd748, -32'd8018, -32'd4690, -32'd10728},
{-32'd2476, 32'd181, -32'd5703, -32'd1790},
{32'd7432, -32'd1928, 32'd3897, 32'd1300},
{32'd1479, 32'd9209, -32'd4230, -32'd2906},
{-32'd13778, -32'd2792, -32'd9091, -32'd14620},
{32'd7683, 32'd316, 32'd4919, 32'd6817},
{32'd4436, 32'd5330, 32'd8175, -32'd7177},
{32'd9874, 32'd498, 32'd1877, -32'd1947},
{-32'd11157, 32'd937, -32'd5696, -32'd7454},
{-32'd6857, 32'd7978, 32'd5504, 32'd1121},
{-32'd4946, -32'd11129, -32'd2724, -32'd6946},
{32'd1141, 32'd31, 32'd11126, -32'd2081},
{32'd4588, -32'd1785, -32'd6289, -32'd9809},
{32'd2733, 32'd1493, -32'd1282, -32'd5777},
{-32'd4033, 32'd1150, -32'd4374, 32'd1056},
{-32'd1722, -32'd9870, -32'd6351, -32'd3737},
{-32'd1680, -32'd14512, 32'd980, 32'd2536},
{-32'd4481, -32'd9436, -32'd2005, -32'd1536},
{-32'd2074, -32'd6762, -32'd5725, -32'd6049},
{-32'd11749, -32'd770, -32'd4478, 32'd4749},
{32'd2298, 32'd897, -32'd10216, 32'd5333},
{-32'd6334, -32'd554, 32'd2113, -32'd767},
{32'd3283, 32'd4311, 32'd6473, -32'd1104},
{-32'd2125, -32'd4716, -32'd4071, 32'd7399},
{32'd4889, 32'd9880, -32'd1006, -32'd3749},
{-32'd4443, -32'd3809, -32'd2412, 32'd872},
{-32'd1845, -32'd4077, 32'd3338, 32'd5362},
{32'd5034, 32'd4985, 32'd2262, -32'd9576},
{32'd7425, -32'd2218, 32'd3340, -32'd4591},
{-32'd2557, -32'd5399, -32'd2081, -32'd2530},
{-32'd1261, 32'd893, -32'd1465, -32'd6369},
{-32'd8520, -32'd5295, -32'd8225, 32'd1132},
{-32'd1277, -32'd3044, -32'd2311, -32'd7584},
{-32'd7711, 32'd8376, 32'd3727, -32'd4858},
{-32'd2745, -32'd4943, 32'd5153, -32'd393},
{32'd6663, 32'd3651, 32'd3162, 32'd1682},
{-32'd4999, 32'd3389, 32'd3823, -32'd1075},
{32'd3886, 32'd2140, 32'd1105, -32'd9923},
{-32'd2665, 32'd748, -32'd4865, 32'd1483},
{-32'd4084, -32'd7689, -32'd68, 32'd4733},
{32'd3328, 32'd6267, 32'd5794, -32'd4347},
{32'd2037, -32'd6971, -32'd3449, -32'd9673},
{-32'd10976, 32'd2209, -32'd6167, 32'd2643},
{32'd3430, 32'd7007, -32'd1919, -32'd2213},
{32'd721, -32'd4994, -32'd4590, 32'd6544},
{-32'd939, 32'd1501, 32'd7412, 32'd4041},
{-32'd4622, -32'd11596, 32'd1324, 32'd445},
{32'd5693, -32'd2292, -32'd2526, -32'd824},
{32'd3251, 32'd2509, -32'd755, -32'd7512},
{-32'd1496, 32'd1658, 32'd349, 32'd2519},
{-32'd11528, -32'd3746, -32'd6574, -32'd476},
{-32'd4463, 32'd12698, 32'd743, -32'd4756},
{32'd9160, -32'd2364, 32'd1459, -32'd5913},
{32'd6417, -32'd3624, 32'd1791, 32'd107},
{-32'd5156, 32'd1035, -32'd4473, -32'd2481},
{32'd1312, -32'd6259, -32'd1889, 32'd5677},
{-32'd5960, 32'd539, 32'd1781, 32'd2963},
{-32'd12242, 32'd4885, -32'd10392, -32'd8999},
{-32'd1798, 32'd4930, 32'd5383, 32'd1936},
{32'd5533, 32'd278, -32'd920, 32'd4944},
{32'd3596, -32'd7874, -32'd1825, 32'd5518},
{-32'd6184, 32'd7034, -32'd608, -32'd4704},
{32'd671, 32'd5448, -32'd3256, -32'd3955},
{32'd917, -32'd3683, -32'd7333, -32'd5735},
{-32'd7949, 32'd5115, 32'd343, 32'd6492},
{-32'd5178, -32'd1747, -32'd1908, -32'd9981},
{-32'd2867, -32'd266, 32'd3164, -32'd5504},
{32'd8673, -32'd5932, -32'd6244, 32'd2596},
{-32'd5790, -32'd5625, 32'd7383, -32'd5677},
{32'd17309, -32'd3322, -32'd2836, 32'd1557},
{32'd7195, 32'd2907, -32'd2060, 32'd322},
{32'd11717, -32'd5590, 32'd8323, -32'd2679},
{-32'd3120, 32'd1155, 32'd9580, 32'd6878},
{32'd5032, 32'd7685, -32'd7184, 32'd2825},
{32'd4625, 32'd968, -32'd1098, 32'd1926},
{32'd7655, 32'd3528, 32'd799, 32'd2881},
{-32'd1663, -32'd1010, -32'd1254, 32'd2207},
{-32'd3083, 32'd1295, 32'd3018, 32'd1318},
{32'd2630, 32'd3365, -32'd3821, -32'd4864},
{-32'd4173, -32'd873, 32'd5464, 32'd3336},
{-32'd2228, 32'd532, -32'd2624, -32'd4354},
{-32'd307, -32'd502, 32'd2062, 32'd3311},
{32'd4636, 32'd5790, 32'd888, 32'd2102},
{32'd1237, -32'd6496, 32'd7664, 32'd10784},
{32'd546, -32'd10951, -32'd10771, -32'd4450},
{-32'd11587, -32'd4665, -32'd6651, 32'd9581},
{-32'd514, 32'd5970, -32'd6722, -32'd4271},
{32'd6305, -32'd4712, -32'd7454, -32'd3414},
{-32'd2761, -32'd613, 32'd3421, -32'd1042},
{-32'd6554, -32'd4944, -32'd6074, 32'd5198},
{32'd9384, 32'd437, -32'd4691, -32'd1234},
{-32'd5514, 32'd2188, 32'd2160, 32'd10364},
{32'd3315, -32'd10459, 32'd1402, -32'd5838},
{-32'd4986, -32'd2737, 32'd2823, 32'd3764},
{32'd11480, 32'd7982, 32'd2543, 32'd2485},
{-32'd2557, -32'd2689, -32'd2387, -32'd6781},
{-32'd2243, -32'd3110, -32'd3342, -32'd1246},
{32'd2827, 32'd7691, -32'd5703, 32'd1584},
{32'd9071, -32'd304, 32'd1382, 32'd1450},
{-32'd4722, -32'd935, -32'd549, -32'd291},
{-32'd7078, -32'd377, -32'd1708, -32'd826},
{32'd4881, 32'd1890, 32'd2192, -32'd3080},
{32'd3708, 32'd3587, 32'd1805, -32'd3404},
{32'd11717, 32'd1592, -32'd3379, 32'd3241},
{-32'd5495, -32'd2822, -32'd5580, -32'd5018},
{32'd526, 32'd2310, 32'd6575, 32'd1081},
{32'd112, 32'd4100, -32'd3840, 32'd2234},
{32'd5081, -32'd4568, 32'd8585, 32'd5385},
{-32'd12703, -32'd2993, 32'd1360, 32'd2355},
{-32'd2836, 32'd7182, -32'd532, -32'd576},
{32'd2157, -32'd2845, 32'd2177, 32'd3902},
{-32'd802, -32'd4418, 32'd2111, -32'd2788},
{-32'd10980, -32'd1713, -32'd4880, -32'd3761},
{32'd3426, -32'd2874, -32'd4068, -32'd1784},
{-32'd583, 32'd3921, -32'd300, 32'd1706},
{32'd10562, 32'd10582, -32'd2059, 32'd1157},
{32'd22841, -32'd5910, 32'd10010, 32'd9376},
{-32'd1583, 32'd4121, 32'd5736, -32'd4656},
{-32'd17418, -32'd2719, -32'd6820, -32'd5636},
{-32'd7410, 32'd2599, 32'd6020, -32'd571},
{32'd3074, -32'd190, -32'd4634, 32'd2265},
{32'd2192, 32'd6189, 32'd5146, 32'd1745},
{-32'd3147, -32'd10241, -32'd5421, -32'd4985},
{-32'd2557, -32'd3388, -32'd1997, 32'd903},
{-32'd439, 32'd3991, -32'd4870, 32'd5175},
{-32'd7568, 32'd563, -32'd3705, -32'd3122},
{32'd4177, 32'd8516, 32'd4246, 32'd5455},
{-32'd4194, -32'd4913, -32'd6202, 32'd1341},
{32'd7421, -32'd6074, 32'd3389, -32'd3480},
{32'd5019, -32'd3442, -32'd1683, 32'd469},
{32'd3272, 32'd7457, -32'd2971, 32'd4591},
{-32'd4336, 32'd1676, 32'd669, -32'd10478},
{32'd1921, -32'd7749, 32'd4593, 32'd11329},
{-32'd4706, -32'd12185, -32'd6602, -32'd5053},
{-32'd1047, 32'd6594, -32'd2812, 32'd8361},
{-32'd8596, -32'd9195, -32'd5934, -32'd2342},
{32'd11324, 32'd2455, 32'd20, -32'd8846},
{-32'd5908, -32'd6861, -32'd12422, -32'd676},
{-32'd5100, -32'd4931, -32'd672, 32'd1720},
{32'd3359, -32'd1039, -32'd6669, -32'd1822},
{32'd4219, -32'd4470, 32'd72, 32'd7209},
{32'd8389, 32'd15978, 32'd4575, -32'd2502},
{32'd581, -32'd4194, -32'd6872, 32'd6137},
{-32'd2741, -32'd4793, -32'd1624, 32'd1508},
{-32'd9497, -32'd2038, -32'd11108, -32'd7655},
{-32'd438, -32'd2829, 32'd2966, 32'd1318},
{-32'd685, -32'd1280, -32'd6145, -32'd4601},
{32'd11509, 32'd3781, 32'd4972, 32'd6094},
{-32'd9583, -32'd3586, 32'd3511, 32'd7539},
{-32'd9374, 32'd5025, -32'd1086, -32'd3043}
},
{{-32'd4095, 32'd6041, 32'd3631, 32'd7014},
{32'd500, -32'd9849, -32'd2391, 32'd100},
{-32'd5780, 32'd1361, -32'd1736, 32'd6473},
{32'd17143, -32'd2327, 32'd2974, -32'd7338},
{-32'd10634, 32'd5960, -32'd3015, 32'd6897},
{32'd6695, -32'd1693, -32'd13720, -32'd9070},
{-32'd3810, 32'd4539, 32'd1095, 32'd4716},
{32'd5025, -32'd13492, -32'd5593, -32'd6790},
{-32'd2747, -32'd105, 32'd2302, 32'd908},
{32'd3112, 32'd6659, 32'd7127, 32'd7628},
{-32'd8463, -32'd3069, -32'd4105, 32'd6934},
{32'd5385, 32'd10003, -32'd3568, -32'd3051},
{32'd9994, 32'd6882, 32'd4638, -32'd3382},
{-32'd497, -32'd11391, -32'd5262, -32'd7756},
{32'd5429, 32'd2176, 32'd1016, -32'd7550},
{32'd1996, 32'd2344, -32'd20528, -32'd8325},
{-32'd4181, 32'd6111, -32'd5163, 32'd3455},
{-32'd5777, -32'd2825, -32'd7931, -32'd2954},
{32'd6912, -32'd3120, -32'd4988, -32'd2165},
{-32'd7008, 32'd6868, 32'd4439, -32'd1701},
{32'd8020, 32'd6864, 32'd4493, 32'd4328},
{32'd3196, -32'd4854, -32'd3311, -32'd6115},
{-32'd6834, -32'd13962, 32'd4456, -32'd12210},
{32'd674, 32'd4316, -32'd9109, -32'd4854},
{32'd480, 32'd11666, 32'd3033, 32'd6841},
{32'd4424, -32'd3673, -32'd266, 32'd9425},
{-32'd4061, 32'd9758, 32'd5919, -32'd3244},
{32'd19717, -32'd7717, 32'd602, -32'd241},
{32'd7409, 32'd6882, 32'd5959, -32'd4232},
{-32'd657, 32'd564, 32'd2123, 32'd287},
{-32'd1548, 32'd5611, -32'd3161, -32'd1324},
{-32'd5133, -32'd6136, -32'd3777, -32'd1814},
{32'd4155, 32'd4953, -32'd6917, 32'd6216},
{32'd4046, 32'd8766, -32'd2484, -32'd6774},
{32'd6977, 32'd13778, 32'd3153, 32'd8441},
{-32'd6209, -32'd8249, -32'd9427, -32'd1388},
{32'd10015, -32'd9014, -32'd11572, 32'd7396},
{32'd7372, -32'd1544, -32'd3998, -32'd6703},
{-32'd1400, 32'd9467, -32'd5093, -32'd1300},
{32'd2992, 32'd9751, -32'd1735, -32'd4774},
{-32'd13152, -32'd214, -32'd4248, 32'd2264},
{32'd1051, 32'd12891, 32'd1890, 32'd4825},
{-32'd9201, 32'd8836, -32'd3887, -32'd13143},
{32'd3876, -32'd775, -32'd6935, -32'd7766},
{-32'd962, -32'd4318, 32'd100, -32'd4773},
{32'd6220, -32'd1611, 32'd422, -32'd9922},
{-32'd7796, -32'd10619, -32'd3448, -32'd7392},
{32'd3362, -32'd5787, -32'd4953, 32'd3603},
{32'd4944, 32'd9688, 32'd2525, 32'd11655},
{-32'd10921, 32'd1517, 32'd9282, 32'd3768},
{-32'd16258, 32'd6924, 32'd2752, 32'd1183},
{32'd13800, 32'd3766, -32'd7448, 32'd2044},
{-32'd5596, -32'd245, -32'd462, 32'd144},
{-32'd8196, 32'd2777, 32'd4526, 32'd1409},
{32'd4175, -32'd1404, 32'd1806, 32'd1342},
{32'd4053, -32'd15290, 32'd2468, 32'd2986},
{32'd9643, 32'd972, 32'd1128, 32'd6769},
{-32'd3859, -32'd6618, -32'd10474, 32'd249},
{-32'd3391, -32'd2476, 32'd4985, -32'd1723},
{-32'd3797, 32'd5457, 32'd6053, -32'd1481},
{-32'd2202, 32'd7796, 32'd6331, 32'd1213},
{32'd15437, -32'd4530, -32'd8086, -32'd8222},
{-32'd10274, -32'd956, -32'd2899, -32'd6114},
{-32'd3941, 32'd3355, 32'd8803, 32'd2137},
{32'd10506, -32'd14, 32'd10369, 32'd6220},
{32'd2522, 32'd14897, 32'd8324, 32'd5366},
{32'd378, -32'd3062, -32'd5096, -32'd2517},
{32'd3693, -32'd291, -32'd1294, 32'd1658},
{32'd5757, -32'd3577, -32'd6754, -32'd5570},
{32'd5084, -32'd1992, 32'd1701, 32'd4027},
{32'd11050, 32'd4364, -32'd1858, -32'd1709},
{32'd10067, -32'd470, -32'd5633, -32'd5550},
{32'd1419, 32'd467, -32'd3225, -32'd2416},
{-32'd4727, 32'd11083, -32'd302, 32'd4579},
{32'd12612, 32'd7857, 32'd10377, 32'd7531},
{-32'd5753, -32'd972, -32'd13819, 32'd613},
{-32'd9520, -32'd4336, -32'd16005, -32'd3126},
{32'd7686, -32'd2903, -32'd8949, 32'd10521},
{32'd2454, 32'd7730, -32'd7216, 32'd6969},
{32'd858, -32'd1138, -32'd8869, 32'd10614},
{32'd3505, 32'd1448, 32'd3476, 32'd4793},
{32'd7855, 32'd4729, -32'd1089, -32'd2385},
{-32'd3377, 32'd338, 32'd7215, -32'd6937},
{-32'd15543, 32'd2503, 32'd11673, 32'd3601},
{-32'd17405, -32'd3888, -32'd4675, -32'd2112},
{-32'd7654, -32'd900, 32'd4755, -32'd488},
{32'd4668, 32'd6293, 32'd11535, -32'd805},
{-32'd3868, -32'd705, -32'd2616, -32'd6871},
{32'd3334, -32'd1670, -32'd996, 32'd5890},
{-32'd2641, -32'd2146, 32'd3064, -32'd2296},
{32'd15128, -32'd898, 32'd2846, -32'd5987},
{-32'd9143, -32'd2650, -32'd4958, 32'd4406},
{32'd6057, 32'd3184, -32'd1341, 32'd2977},
{32'd8379, 32'd6076, 32'd5132, 32'd3280},
{32'd2412, -32'd5287, 32'd1415, -32'd1900},
{32'd1564, -32'd11704, 32'd4409, 32'd10720},
{32'd1898, 32'd11458, -32'd10032, 32'd3109},
{-32'd12224, -32'd4151, -32'd8178, 32'd3381},
{32'd9348, 32'd7981, 32'd1839, 32'd5569},
{-32'd328, 32'd4207, -32'd383, -32'd2737},
{-32'd5156, -32'd1745, -32'd14160, -32'd5190},
{-32'd6760, -32'd2795, 32'd10836, 32'd7281},
{-32'd1066, -32'd1411, -32'd5351, -32'd5652},
{32'd5923, 32'd16574, -32'd2772, 32'd3404},
{-32'd328, 32'd9898, -32'd2334, -32'd456},
{32'd3730, 32'd3401, -32'd6177, 32'd2276},
{32'd5781, -32'd5742, -32'd1781, 32'd4092},
{-32'd11428, -32'd1497, 32'd6204, -32'd7315},
{-32'd4111, 32'd6978, -32'd1518, 32'd5626},
{-32'd14486, -32'd4025, 32'd871, 32'd6957},
{-32'd11993, 32'd9022, 32'd321, -32'd1455},
{-32'd4679, 32'd11296, 32'd1151, -32'd3823},
{32'd5604, -32'd1198, -32'd2512, 32'd2775},
{-32'd1612, 32'd2875, 32'd9945, 32'd1500},
{-32'd10898, -32'd5081, 32'd5198, -32'd2389},
{-32'd12306, -32'd1114, 32'd3075, 32'd678},
{-32'd5147, -32'd5389, 32'd10108, 32'd6836},
{-32'd6358, -32'd6847, 32'd301, -32'd67},
{32'd8945, 32'd2232, 32'd768, -32'd18182},
{32'd9470, 32'd7186, -32'd5203, 32'd8161},
{32'd1650, 32'd346, -32'd10973, -32'd6739},
{-32'd1547, 32'd196, -32'd6921, 32'd1772},
{32'd6541, 32'd2511, -32'd6319, -32'd3511},
{-32'd1204, -32'd13055, 32'd982, -32'd3368},
{32'd8576, -32'd4605, 32'd4670, 32'd6162},
{32'd4192, -32'd2179, 32'd12446, -32'd2914},
{-32'd12895, -32'd8995, -32'd6114, -32'd677},
{32'd5572, -32'd3219, 32'd1921, -32'd3091},
{-32'd15322, -32'd13165, 32'd1722, -32'd4887},
{32'd6053, 32'd9084, 32'd1252, 32'd7972},
{-32'd14411, 32'd6726, 32'd8500, 32'd734},
{-32'd6853, -32'd6468, -32'd1163, -32'd2599},
{-32'd3243, -32'd4117, -32'd1542, -32'd515},
{32'd6801, 32'd9050, -32'd2552, -32'd6551},
{32'd21052, 32'd864, -32'd3044, -32'd4724},
{-32'd2073, 32'd252, -32'd6527, 32'd8941},
{32'd8947, 32'd1501, 32'd1291, -32'd7353},
{-32'd2722, -32'd2614, -32'd2919, 32'd5342},
{32'd5334, -32'd7114, 32'd9474, -32'd2633},
{32'd4611, -32'd6370, -32'd3101, -32'd1119},
{32'd12116, 32'd7745, 32'd10186, 32'd7361},
{-32'd628, 32'd4821, -32'd12827, -32'd7112},
{-32'd13777, -32'd8511, 32'd8208, -32'd5269},
{32'd8408, -32'd3075, 32'd6706, 32'd1980},
{32'd1597, 32'd4804, -32'd127, 32'd3769},
{-32'd4736, 32'd12142, 32'd3076, -32'd2388},
{-32'd7630, 32'd4666, -32'd6046, 32'd3513},
{-32'd20351, 32'd2097, -32'd7668, -32'd2969},
{32'd5757, 32'd4369, 32'd709, -32'd8110},
{32'd7900, -32'd8444, -32'd449, -32'd14},
{32'd3306, -32'd8071, -32'd6722, -32'd3280},
{-32'd4516, 32'd4153, 32'd3622, -32'd307},
{-32'd13293, 32'd47, -32'd7404, -32'd97},
{-32'd6463, 32'd5886, 32'd1469, 32'd12433},
{-32'd1199, -32'd1207, 32'd6190, -32'd9286},
{32'd2293, -32'd15365, -32'd3674, -32'd4796},
{-32'd1002, 32'd9578, -32'd511, 32'd6438},
{32'd8728, -32'd8416, 32'd15599, 32'd8285},
{-32'd4768, 32'd5083, 32'd1721, -32'd5147},
{32'd6423, 32'd3917, -32'd564, 32'd5014},
{-32'd7010, -32'd10065, -32'd11374, 32'd10157},
{32'd5916, -32'd8875, -32'd4513, -32'd5270},
{-32'd8344, -32'd797, -32'd7637, -32'd15487},
{32'd8962, 32'd9281, 32'd7434, -32'd3847},
{-32'd8861, 32'd11926, 32'd3779, 32'd1182},
{-32'd3385, 32'd5810, 32'd2276, 32'd1250},
{-32'd3545, 32'd6301, 32'd9501, 32'd8882},
{-32'd3618, -32'd2031, -32'd3125, -32'd4221},
{-32'd262, -32'd1094, -32'd761, -32'd7060},
{32'd4520, -32'd3686, -32'd5142, -32'd5517},
{32'd5660, -32'd9477, 32'd2490, -32'd4584},
{32'd9419, 32'd6253, 32'd10419, -32'd3280},
{32'd6551, 32'd6365, 32'd3083, 32'd6306},
{32'd3652, -32'd8590, 32'd172, 32'd1583},
{32'd9992, 32'd10866, 32'd11235, -32'd2621},
{-32'd3810, -32'd5303, -32'd15669, 32'd8689},
{32'd3240, -32'd10711, 32'd13309, -32'd4585},
{32'd5748, 32'd2929, -32'd8406, -32'd9060},
{-32'd10425, -32'd1400, -32'd3163, -32'd3973},
{32'd70, -32'd12742, -32'd70, -32'd7042},
{-32'd12936, 32'd12184, 32'd5822, -32'd2278},
{-32'd3933, -32'd6103, -32'd6920, -32'd2891},
{-32'd3695, -32'd2587, -32'd10269, -32'd2673},
{32'd3338, 32'd2880, -32'd962, -32'd10839},
{-32'd5314, -32'd769, -32'd1176, 32'd4259},
{-32'd4545, -32'd3683, 32'd5152, 32'd7360},
{32'd5478, 32'd2099, 32'd10703, -32'd1725},
{32'd6786, 32'd4579, 32'd2630, -32'd4036},
{-32'd4528, 32'd1585, -32'd4323, -32'd2636},
{-32'd1039, -32'd15411, -32'd4222, -32'd322},
{32'd5430, 32'd1376, -32'd6520, -32'd6599},
{32'd6435, 32'd4015, -32'd11949, -32'd1463},
{-32'd8361, 32'd6389, -32'd2946, -32'd563},
{32'd4278, 32'd11165, -32'd3013, -32'd1373},
{32'd989, -32'd898, -32'd3874, 32'd2879},
{32'd3061, 32'd3532, 32'd2375, -32'd1909},
{-32'd2916, 32'd1634, -32'd3254, -32'd144},
{32'd3049, 32'd2080, -32'd4376, 32'd3016},
{32'd3979, -32'd11658, -32'd3181, 32'd634},
{-32'd2502, -32'd3533, -32'd12052, -32'd3987},
{-32'd1155, -32'd15660, -32'd7267, -32'd5989},
{32'd846, 32'd9070, -32'd442, -32'd3666},
{32'd10756, 32'd10954, -32'd324, -32'd1957},
{32'd4841, 32'd539, -32'd6520, -32'd981},
{32'd8830, -32'd3666, -32'd8743, -32'd4003},
{32'd11699, -32'd5817, 32'd5246, 32'd10791},
{-32'd1168, 32'd3222, -32'd1390, 32'd4734},
{32'd194, -32'd8926, -32'd3529, -32'd8352},
{32'd8082, -32'd12284, -32'd14342, 32'd2128},
{-32'd7487, 32'd5858, -32'd4304, 32'd109},
{32'd11665, 32'd5826, -32'd3824, 32'd2964},
{-32'd4430, -32'd2045, -32'd6093, 32'd2595},
{-32'd3348, 32'd2640, 32'd9686, 32'd5952},
{-32'd536, 32'd5646, -32'd1835, -32'd997},
{-32'd6063, 32'd1916, 32'd4598, -32'd13711},
{-32'd3449, 32'd9358, -32'd5235, -32'd6664},
{32'd3578, 32'd442, 32'd11266, -32'd9350},
{-32'd2143, 32'd3072, 32'd690, -32'd312},
{32'd4259, 32'd6470, 32'd5296, 32'd1430},
{32'd514, 32'd4158, -32'd4202, -32'd4635},
{-32'd4195, 32'd820, -32'd5144, -32'd6108},
{-32'd17863, 32'd1108, 32'd6976, 32'd5063},
{-32'd1131, 32'd6361, 32'd1370, 32'd4353},
{-32'd2428, 32'd1204, 32'd4086, -32'd593},
{32'd1250, -32'd2095, -32'd310, 32'd5330},
{32'd14338, 32'd524, -32'd7001, 32'd1102},
{-32'd6262, -32'd3606, -32'd1150, -32'd554},
{32'd4184, 32'd2215, -32'd4698, -32'd3247},
{32'd5714, -32'd3861, -32'd4218, -32'd12049},
{32'd2860, 32'd909, 32'd5786, 32'd1463},
{-32'd9373, 32'd14517, 32'd8158, 32'd8311},
{-32'd9236, 32'd2951, 32'd7903, -32'd1937},
{32'd8000, 32'd2316, -32'd697, 32'd11007},
{-32'd14886, -32'd8615, 32'd485, 32'd4151},
{-32'd2712, -32'd9066, -32'd2146, -32'd8252},
{-32'd10176, -32'd16973, 32'd6737, -32'd5262},
{-32'd8198, -32'd9967, -32'd2799, 32'd4714},
{32'd8939, -32'd684, -32'd5237, -32'd4775},
{-32'd338, 32'd10156, 32'd8666, -32'd86},
{-32'd5130, -32'd12603, -32'd13598, 32'd1263},
{-32'd1310, 32'd9366, -32'd525, 32'd872},
{-32'd6298, -32'd5929, -32'd3956, 32'd5526},
{32'd418, -32'd15415, -32'd3215, -32'd7229},
{32'd8196, 32'd3271, 32'd10736, -32'd910},
{32'd8211, 32'd5338, 32'd6231, 32'd13468},
{32'd2203, -32'd5191, -32'd3738, -32'd1028},
{-32'd1065, -32'd5240, -32'd762, -32'd6156},
{-32'd2759, -32'd3520, 32'd950, 32'd5172},
{32'd7401, -32'd11601, -32'd10848, 32'd2669},
{-32'd1384, -32'd3907, 32'd2117, -32'd5094},
{32'd672, -32'd3287, 32'd7949, 32'd3210},
{32'd714, -32'd4187, -32'd3860, 32'd10660},
{-32'd6820, 32'd6304, -32'd4982, 32'd222},
{32'd3424, 32'd7992, 32'd997, -32'd766},
{-32'd6551, 32'd4990, 32'd2694, -32'd9989},
{32'd7331, 32'd11780, -32'd375, -32'd5324},
{-32'd10521, 32'd6348, 32'd8441, 32'd962},
{32'd14375, 32'd5046, 32'd3483, -32'd4592},
{-32'd4087, -32'd2376, 32'd3942, -32'd4381},
{32'd3014, 32'd2822, 32'd1743, -32'd5573},
{32'd2615, -32'd5724, 32'd9471, -32'd5404},
{-32'd13967, 32'd142, -32'd9808, 32'd1221},
{-32'd10068, -32'd967, -32'd4600, 32'd109},
{32'd8208, 32'd936, -32'd10228, -32'd4103},
{32'd1339, 32'd5240, 32'd1510, 32'd2304},
{-32'd736, -32'd6217, -32'd1657, 32'd2719},
{-32'd4106, -32'd1950, -32'd1611, 32'd69},
{-32'd4063, -32'd2103, 32'd2612, 32'd7976},
{-32'd5780, -32'd1801, 32'd1482, 32'd2248},
{-32'd4813, -32'd7301, 32'd873, 32'd2681},
{-32'd1791, -32'd4028, 32'd3095, 32'd5911},
{32'd906, 32'd2502, 32'd5911, 32'd7141},
{-32'd2603, 32'd1829, -32'd4148, -32'd1543},
{-32'd10862, 32'd4698, -32'd1838, -32'd2183},
{-32'd11552, 32'd7137, 32'd2579, 32'd3369},
{-32'd8336, -32'd1590, -32'd1145, 32'd3051},
{32'd3741, 32'd12275, 32'd6443, 32'd10326},
{-32'd2133, 32'd6115, -32'd7928, -32'd7547},
{-32'd5237, -32'd8971, -32'd9325, -32'd4557},
{32'd4758, -32'd7899, -32'd8261, 32'd1433},
{32'd1269, 32'd3893, -32'd6221, -32'd962},
{-32'd7603, -32'd708, 32'd9561, 32'd3416},
{32'd4422, -32'd8879, 32'd5320, 32'd767},
{32'd9637, 32'd4873, 32'd137, 32'd6309},
{-32'd4495, 32'd7392, 32'd6610, -32'd588},
{-32'd8447, -32'd14048, -32'd4145, -32'd12601},
{-32'd202, -32'd4831, 32'd16470, 32'd1236},
{-32'd9584, -32'd7405, -32'd8759, -32'd2252},
{-32'd3752, -32'd471, -32'd9947, -32'd5918},
{-32'd20192, -32'd1566, -32'd11319, 32'd1422},
{-32'd3540, 32'd3637, 32'd2626, 32'd2795},
{32'd11257, 32'd5180, 32'd3287, 32'd188},
{-32'd2095, -32'd7616, 32'd4167, 32'd674},
{-32'd8111, -32'd5410, -32'd7166, 32'd503},
{32'd5600, -32'd11862, -32'd998, -32'd8839},
{-32'd2899, -32'd3887, -32'd4341, -32'd5946},
{32'd3095, 32'd4634, 32'd5440, 32'd517},
{32'd4844, 32'd4307, 32'd4802, -32'd764},
{32'd10996, 32'd7769, -32'd3835, -32'd2045},
{-32'd14985, 32'd176, -32'd11153, -32'd524}
},
{{32'd609, -32'd2491, 32'd2213, -32'd1461},
{-32'd10916, -32'd11032, -32'd8482, 32'd2607},
{-32'd5260, 32'd1317, -32'd11217, 32'd11348},
{32'd390, 32'd13025, 32'd614, 32'd10143},
{32'd10023, 32'd7683, -32'd1440, 32'd5481},
{-32'd7005, -32'd5564, 32'd12997, -32'd7647},
{32'd547, -32'd4668, 32'd6218, 32'd1637},
{-32'd5726, -32'd5171, -32'd10991, -32'd8874},
{32'd6573, 32'd534, -32'd955, 32'd3081},
{32'd15269, 32'd6826, 32'd5271, 32'd5123},
{-32'd1904, -32'd8398, -32'd3749, 32'd1624},
{-32'd388, -32'd1084, 32'd1854, 32'd1613},
{-32'd4207, 32'd5266, 32'd2578, -32'd4636},
{-32'd5480, -32'd2030, -32'd4678, 32'd4262},
{32'd3320, 32'd12458, -32'd5548, 32'd1025},
{-32'd2350, -32'd7098, 32'd10791, -32'd2113},
{-32'd635, 32'd18378, 32'd1410, 32'd16970},
{-32'd2921, -32'd6391, 32'd3440, -32'd15857},
{-32'd3586, -32'd2203, 32'd1265, 32'd9402},
{32'd2675, 32'd4826, -32'd3923, 32'd1253},
{32'd3627, 32'd8673, 32'd5124, 32'd2090},
{-32'd14610, -32'd10574, -32'd6836, -32'd9225},
{-32'd270, -32'd9347, -32'd150, -32'd4580},
{-32'd5596, 32'd11250, -32'd7328, -32'd3067},
{32'd8665, -32'd4381, 32'd5376, 32'd2989},
{32'd7094, 32'd17419, 32'd11070, 32'd6412},
{32'd528, -32'd9134, 32'd1164, -32'd3284},
{-32'd1895, -32'd445, 32'd1605, 32'd4964},
{-32'd5188, -32'd418, -32'd263, 32'd4917},
{32'd8086, -32'd17499, 32'd3319, -32'd13009},
{-32'd7480, 32'd5314, 32'd11952, 32'd496},
{-32'd8953, -32'd5522, -32'd5750, -32'd6624},
{32'd5664, -32'd806, -32'd4842, 32'd1051},
{-32'd1988, -32'd3422, -32'd2190, -32'd4588},
{32'd9127, 32'd5619, 32'd12987, -32'd3573},
{32'd3000, 32'd2883, -32'd3179, 32'd9557},
{-32'd1599, 32'd7883, -32'd8546, 32'd2512},
{32'd10290, 32'd4453, 32'd3645, 32'd5408},
{32'd4662, 32'd190, -32'd12418, -32'd4964},
{-32'd4729, -32'd3294, -32'd15908, -32'd7987},
{32'd1729, 32'd1730, -32'd9910, 32'd1532},
{32'd6558, -32'd1378, -32'd1562, 32'd1009},
{-32'd5840, -32'd576, 32'd4290, -32'd569},
{-32'd6042, -32'd6465, 32'd4604, -32'd1568},
{32'd2321, -32'd9162, -32'd8402, -32'd4791},
{-32'd2891, -32'd2061, 32'd11234, -32'd5748},
{-32'd7415, -32'd14241, -32'd729, 32'd8201},
{32'd2629, 32'd4312, -32'd6613, 32'd462},
{32'd1624, 32'd9552, 32'd13172, -32'd5407},
{32'd496, 32'd870, -32'd5005, -32'd204},
{-32'd6235, -32'd2168, -32'd9487, 32'd431},
{-32'd715, 32'd8820, 32'd2892, 32'd8324},
{-32'd8347, -32'd4982, 32'd1384, 32'd508},
{-32'd4213, -32'd712, -32'd6248, -32'd2089},
{32'd3065, 32'd4928, 32'd9918, 32'd1992},
{-32'd12329, -32'd1065, -32'd11830, -32'd636},
{32'd4726, 32'd1692, -32'd7335, 32'd14748},
{32'd6654, -32'd12023, 32'd853, -32'd2572},
{-32'd8788, -32'd11322, -32'd7529, -32'd6897},
{32'd2684, -32'd7653, 32'd1761, -32'd1528},
{32'd496, 32'd6661, 32'd7670, 32'd1237},
{-32'd9494, 32'd6339, -32'd8765, 32'd6718},
{32'd4323, 32'd5897, -32'd6133, -32'd971},
{32'd11862, -32'd1306, -32'd7037, 32'd5882},
{32'd7114, 32'd1450, -32'd1581, 32'd2911},
{32'd5953, 32'd3619, 32'd6838, -32'd40},
{32'd2961, 32'd3834, 32'd11453, -32'd5982},
{-32'd4427, 32'd1430, -32'd420, -32'd4203},
{32'd8112, -32'd1063, -32'd379, -32'd703},
{32'd2962, 32'd4584, 32'd249, -32'd5679},
{32'd797, -32'd5626, -32'd7179, -32'd3187},
{-32'd2126, -32'd505, -32'd11795, -32'd3342},
{-32'd1173, -32'd3323, -32'd4467, 32'd2756},
{-32'd2445, -32'd2991, -32'd14554, -32'd1345},
{32'd1983, 32'd5443, 32'd4617, 32'd1194},
{32'd2013, -32'd6429, 32'd3804, -32'd3627},
{-32'd4196, -32'd16612, -32'd16377, 32'd3098},
{-32'd1781, 32'd5158, 32'd3433, 32'd6838},
{-32'd4654, 32'd8524, 32'd10327, 32'd4254},
{32'd3227, 32'd4583, -32'd7092, 32'd4580},
{32'd7582, -32'd13356, 32'd7022, 32'd5958},
{-32'd2507, -32'd5044, -32'd4468, 32'd4289},
{-32'd5434, -32'd2387, -32'd5499, 32'd2251},
{32'd1655, -32'd1787, 32'd4764, 32'd601},
{-32'd3132, -32'd10269, -32'd278, -32'd6886},
{32'd7943, 32'd4447, -32'd669, 32'd380},
{32'd5790, 32'd1118, -32'd4160, -32'd3534},
{-32'd731, -32'd9206, -32'd4496, -32'd4687},
{32'd9534, -32'd95, -32'd2284, -32'd7785},
{-32'd5401, 32'd3769, -32'd10019, -32'd2495},
{32'd2408, -32'd6674, -32'd1504, 32'd8875},
{32'd8838, -32'd9749, -32'd4448, 32'd8974},
{32'd1137, 32'd9951, 32'd9858, -32'd1393},
{32'd235, 32'd4591, 32'd12563, 32'd5963},
{32'd1857, 32'd235, -32'd10314, 32'd7116},
{-32'd5575, -32'd2631, 32'd5048, 32'd516},
{32'd4581, 32'd11086, 32'd3910, 32'd8117},
{32'd4965, 32'd7632, 32'd201, 32'd6868},
{-32'd3693, -32'd7825, -32'd3054, -32'd7668},
{32'd10707, 32'd9982, 32'd12454, -32'd2125},
{-32'd462, -32'd1996, 32'd2467, -32'd12388},
{-32'd8657, -32'd9583, 32'd570, -32'd3915},
{32'd4214, -32'd2816, 32'd3462, 32'd1610},
{32'd3791, 32'd2295, 32'd5400, 32'd5087},
{32'd519, 32'd6214, 32'd4529, 32'd5004},
{32'd2545, 32'd3373, 32'd2648, -32'd5485},
{32'd1255, -32'd3382, -32'd3500, -32'd1482},
{32'd1408, 32'd3454, -32'd2684, 32'd12314},
{32'd1262, 32'd10455, 32'd4375, -32'd3863},
{-32'd2840, 32'd1481, -32'd10799, 32'd1973},
{32'd421, -32'd2518, 32'd53, 32'd7462},
{-32'd1483, -32'd9787, -32'd6387, -32'd3925},
{-32'd382, 32'd2514, -32'd3595, 32'd5539},
{32'd3296, 32'd1048, -32'd1152, 32'd4873},
{-32'd573, -32'd5473, -32'd5001, -32'd1193},
{32'd3999, -32'd4494, 32'd169, -32'd9066},
{32'd3806, 32'd9156, 32'd6981, -32'd6344},
{-32'd14625, -32'd18674, -32'd4348, -32'd10259},
{32'd1629, 32'd1001, -32'd4928, 32'd490},
{32'd5739, 32'd7112, 32'd2157, 32'd3153},
{32'd6058, 32'd10924, 32'd5396, -32'd1014},
{-32'd874, 32'd17421, 32'd124, 32'd9728},
{32'd4816, -32'd9141, 32'd4818, -32'd3163},
{-32'd1795, 32'd3352, -32'd6825, 32'd2103},
{-32'd1961, -32'd5318, -32'd3096, 32'd2528},
{32'd2053, -32'd1384, -32'd1575, 32'd1759},
{32'd1705, 32'd2691, -32'd1842, -32'd9150},
{-32'd2071, 32'd2344, -32'd10445, -32'd4304},
{-32'd2423, -32'd10154, -32'd9587, 32'd6363},
{-32'd6693, 32'd6540, -32'd2856, 32'd1400},
{-32'd909, 32'd228, -32'd6157, 32'd1965},
{-32'd3700, -32'd11326, -32'd6137, -32'd8163},
{-32'd1679, -32'd2376, 32'd5498, -32'd10228},
{32'd1346, -32'd4540, -32'd11372, -32'd4673},
{32'd2863, 32'd3673, 32'd3047, 32'd777},
{-32'd2966, 32'd146, -32'd6545, -32'd4128},
{-32'd5779, -32'd7554, -32'd3949, 32'd5525},
{-32'd13894, -32'd245, 32'd3169, 32'd976},
{-32'd4999, 32'd3383, 32'd5205, -32'd2131},
{-32'd641, 32'd938, -32'd5294, 32'd7251},
{32'd5138, 32'd258, -32'd3413, 32'd10404},
{-32'd12215, 32'd5811, -32'd11516, 32'd6698},
{32'd14318, -32'd5849, 32'd3856, 32'd8343},
{-32'd8311, -32'd6145, -32'd10164, 32'd5356},
{32'd7337, 32'd21014, -32'd1782, 32'd80},
{32'd7270, -32'd1502, -32'd3290, 32'd7759},
{-32'd5494, 32'd1290, -32'd5686, -32'd2837},
{32'd7383, -32'd2089, -32'd11973, -32'd7656},
{32'd11549, 32'd447, -32'd2688, -32'd3563},
{-32'd3973, -32'd14929, -32'd8790, -32'd5594},
{-32'd9356, 32'd7112, -32'd386, 32'd454},
{-32'd9973, 32'd5947, 32'd5282, -32'd3698},
{-32'd5698, -32'd4607, -32'd340, -32'd494},
{32'd3466, -32'd7794, 32'd3185, -32'd3053},
{-32'd8320, -32'd20006, -32'd374, -32'd6435},
{32'd3964, 32'd1510, 32'd3588, 32'd2736},
{32'd2008, 32'd5222, -32'd1541, 32'd12898},
{32'd5458, 32'd4963, -32'd1547, -32'd12300},
{32'd2747, -32'd7794, 32'd1119, -32'd5902},
{32'd4187, -32'd3942, -32'd999, 32'd3091},
{-32'd1773, -32'd5271, -32'd1971, 32'd11060},
{32'd119, 32'd7499, -32'd2800, 32'd5398},
{32'd4332, -32'd1875, -32'd1172, -32'd9270},
{-32'd3497, 32'd3801, 32'd629, -32'd1195},
{32'd7055, -32'd1717, -32'd3049, -32'd1321},
{32'd7376, -32'd13537, -32'd8252, -32'd71},
{32'd11208, -32'd1479, 32'd16305, -32'd11815},
{-32'd6347, -32'd10950, -32'd7182, 32'd6192},
{-32'd7145, -32'd1468, 32'd2646, 32'd1220},
{-32'd251, 32'd6855, -32'd2777, -32'd872},
{-32'd7810, 32'd8900, -32'd6401, -32'd3190},
{-32'd5110, -32'd8230, -32'd793, -32'd6249},
{32'd9908, -32'd186, 32'd10876, -32'd2012},
{-32'd2573, 32'd5092, -32'd11058, 32'd904},
{32'd2188, 32'd13568, 32'd1502, 32'd3740},
{32'd3755, -32'd6902, -32'd8666, -32'd2020},
{32'd13006, 32'd5864, -32'd248, -32'd435},
{-32'd1990, -32'd1947, 32'd6194, 32'd89},
{32'd6262, -32'd1817, -32'd928, 32'd5947},
{-32'd1409, 32'd62, -32'd9030, -32'd1911},
{-32'd5640, 32'd9198, -32'd5691, 32'd3314},
{32'd1390, -32'd10746, -32'd5083, 32'd3774},
{-32'd1330, -32'd12438, 32'd5062, -32'd3182},
{32'd811, 32'd1169, -32'd3849, -32'd7996},
{32'd2700, -32'd485, -32'd2609, -32'd4237},
{32'd12161, -32'd3106, 32'd4788, -32'd7135},
{32'd3425, 32'd3963, 32'd1444, -32'd3777},
{-32'd10174, -32'd7061, 32'd3708, 32'd3250},
{32'd6893, -32'd10305, 32'd1174, -32'd10988},
{-32'd2820, -32'd1354, 32'd641, -32'd1787},
{32'd2169, -32'd1238, 32'd6769, -32'd4092},
{-32'd4763, -32'd1022, -32'd7873, -32'd1683},
{32'd10587, 32'd2466, -32'd1689, -32'd1054},
{-32'd1953, -32'd2474, -32'd4081, -32'd10688},
{32'd7923, -32'd7353, -32'd3437, 32'd1585},
{32'd2771, -32'd507, 32'd1790, 32'd11272},
{32'd4923, 32'd6154, -32'd136, 32'd9595},
{-32'd1766, 32'd7253, -32'd2489, 32'd4091},
{-32'd602, 32'd3928, -32'd3530, 32'd8514},
{32'd4729, -32'd1253, 32'd13681, 32'd5877},
{-32'd11104, -32'd7764, -32'd2704, 32'd821},
{32'd4523, 32'd4292, -32'd1243, 32'd2734},
{32'd4416, -32'd331, 32'd1163, -32'd3445},
{32'd3385, 32'd3579, -32'd641, 32'd13836},
{32'd4722, -32'd8557, -32'd2522, -32'd3227},
{-32'd5653, 32'd238, -32'd11883, -32'd10930},
{-32'd5241, 32'd2368, 32'd3079, 32'd5226},
{32'd6551, 32'd1343, -32'd10607, -32'd8075},
{-32'd7904, 32'd5318, -32'd1425, 32'd15611},
{32'd3754, 32'd6072, 32'd14287, -32'd3352},
{-32'd1220, -32'd7515, -32'd903, -32'd3195},
{32'd6486, 32'd3602, 32'd7537, -32'd1530},
{-32'd6697, -32'd3744, -32'd2388, -32'd607},
{32'd3233, 32'd3230, 32'd4434, -32'd1846},
{-32'd3069, -32'd3551, -32'd5797, -32'd2227},
{-32'd5255, 32'd7971, -32'd3824, -32'd1595},
{-32'd1375, -32'd2657, -32'd2212, 32'd3349},
{32'd7959, 32'd6324, -32'd3297, -32'd5876},
{-32'd1854, 32'd11473, -32'd5455, 32'd10490},
{32'd10697, 32'd2264, -32'd4686, -32'd863},
{-32'd1819, -32'd7899, 32'd7039, -32'd499},
{32'd4209, 32'd15539, 32'd1822, 32'd10532},
{32'd540, 32'd627, 32'd6076, 32'd2123},
{32'd4563, -32'd12510, 32'd10530, 32'd613},
{32'd2956, -32'd1277, 32'd10259, 32'd3538},
{-32'd6426, -32'd9437, -32'd5371, -32'd678},
{-32'd4087, -32'd890, 32'd5823, 32'd1521},
{32'd13430, -32'd7463, -32'd5889, -32'd14627},
{-32'd248, -32'd3196, 32'd904, 32'd5426},
{32'd9386, 32'd1011, 32'd4469, 32'd13288},
{-32'd7574, -32'd9182, -32'd12394, -32'd2673},
{-32'd5619, 32'd4121, -32'd8167, 32'd3812},
{32'd2957, 32'd12247, 32'd5342, 32'd12395},
{32'd6129, -32'd279, -32'd1350, 32'd3495},
{-32'd9219, -32'd12145, 32'd1390, -32'd7592},
{32'd2580, -32'd14547, 32'd3122, -32'd18559},
{-32'd7910, -32'd17116, -32'd19299, -32'd5928},
{32'd37, 32'd2032, -32'd1573, -32'd3039},
{-32'd3786, 32'd7841, 32'd15925, 32'd8400},
{-32'd5706, 32'd11181, -32'd6301, 32'd7545},
{32'd7825, -32'd4629, 32'd216, 32'd4393},
{32'd913, 32'd3791, 32'd5196, 32'd4281},
{-32'd13695, 32'd7915, -32'd1665, 32'd1291},
{32'd5275, -32'd2709, -32'd604, 32'd3249},
{32'd13454, -32'd1406, 32'd6360, 32'd2351},
{32'd10752, 32'd11875, -32'd10184, 32'd4550},
{-32'd11197, 32'd1366, 32'd137, -32'd1561},
{32'd3880, -32'd4967, 32'd5512, 32'd2676},
{-32'd6010, 32'd4053, 32'd9393, 32'd3433},
{32'd3750, 32'd6133, 32'd1100, -32'd4652},
{32'd300, -32'd9200, -32'd10521, 32'd4905},
{-32'd1796, 32'd2091, 32'd4492, 32'd2100},
{32'd1084, 32'd3273, 32'd14184, 32'd3702},
{32'd3421, 32'd7214, 32'd10675, 32'd2655},
{-32'd2296, -32'd3967, -32'd7414, -32'd2147},
{-32'd1949, -32'd484, 32'd6487, 32'd984},
{32'd2642, -32'd209, -32'd3710, -32'd1984},
{32'd2315, 32'd3622, 32'd9549, -32'd1304},
{-32'd1434, 32'd1717, -32'd5263, -32'd1240},
{-32'd7017, -32'd7081, -32'd2597, 32'd3154},
{-32'd27, -32'd4359, -32'd1798, -32'd6796},
{32'd7123, 32'd6127, 32'd2611, -32'd6564},
{-32'd3597, 32'd4246, 32'd6213, 32'd6229},
{-32'd2948, 32'd3093, 32'd1962, 32'd8869},
{32'd926, -32'd5264, 32'd1577, 32'd3246},
{-32'd6272, -32'd10405, -32'd9357, 32'd1119},
{-32'd2727, 32'd4998, -32'd4507, -32'd10769},
{32'd11086, 32'd3134, 32'd734, 32'd1874},
{-32'd4533, -32'd3291, 32'd4763, -32'd3336},
{-32'd3060, -32'd418, -32'd18621, 32'd11482},
{-32'd10271, 32'd632, 32'd3047, -32'd2753},
{32'd7966, 32'd2835, -32'd1316, -32'd1531},
{-32'd6680, -32'd2388, -32'd11925, -32'd7367},
{32'd2573, 32'd7241, 32'd10020, -32'd4126},
{-32'd3971, -32'd1066, 32'd2126, 32'd3542},
{-32'd4255, -32'd11122, 32'd107, -32'd4362},
{32'd14010, 32'd5847, 32'd3795, 32'd2806},
{32'd154, 32'd3654, 32'd10518, -32'd4219},
{-32'd8985, 32'd5180, 32'd4423, -32'd4589},
{-32'd7293, 32'd2857, 32'd4520, -32'd4581},
{32'd3522, 32'd5496, 32'd7620, 32'd5301},
{32'd5980, -32'd532, -32'd1195, 32'd813},
{-32'd8342, 32'd3624, 32'd3970, 32'd10568},
{-32'd2925, 32'd2957, -32'd3251, -32'd2908},
{32'd9177, 32'd3504, -32'd749, 32'd586},
{-32'd9253, 32'd904, -32'd10495, 32'd7941},
{-32'd5730, -32'd1450, 32'd8298, -32'd2381},
{32'd2048, -32'd1833, -32'd1061, 32'd2250},
{-32'd2163, 32'd13136, 32'd15268, 32'd9804},
{-32'd6249, 32'd4129, 32'd1355, 32'd660},
{-32'd4374, 32'd375, 32'd2743, -32'd832},
{-32'd5532, 32'd3472, -32'd6412, 32'd5585},
{-32'd3167, 32'd2017, -32'd5252, 32'd6583},
{-32'd1987, -32'd10086, -32'd5270, -32'd5914},
{-32'd2593, 32'd9781, -32'd8780, -32'd3988},
{32'd378, 32'd8514, 32'd1100, -32'd5461},
{-32'd7782, -32'd1298, -32'd278, 32'd3671},
{-32'd725, 32'd4651, 32'd13013, -32'd6884},
{32'd12316, 32'd9592, 32'd450, -32'd4371},
{32'd4033, 32'd3684, -32'd1081, -32'd5917}
},
{{32'd7051, 32'd9662, 32'd2448, -32'd4042},
{-32'd3830, -32'd865, 32'd137, -32'd2154},
{32'd3781, -32'd397, 32'd2812, 32'd5428},
{32'd3227, 32'd4318, 32'd6873, -32'd2111},
{-32'd3152, 32'd1109, -32'd1530, -32'd3741},
{-32'd6561, -32'd8730, 32'd588, -32'd2662},
{32'd6793, 32'd7197, 32'd1968, 32'd4046},
{32'd2371, -32'd5837, -32'd8021, 32'd214},
{-32'd2873, 32'd2523, -32'd6231, -32'd5301},
{32'd13580, 32'd3932, 32'd3357, 32'd7161},
{-32'd9399, 32'd875, -32'd1281, 32'd2006},
{32'd125, -32'd4700, 32'd1530, 32'd1287},
{32'd5347, 32'd3886, -32'd2138, -32'd4092},
{32'd3481, 32'd3055, -32'd4838, -32'd5549},
{32'd1947, 32'd3036, 32'd1120, -32'd4614},
{-32'd756, -32'd1799, 32'd1538, -32'd7691},
{-32'd2732, -32'd1911, -32'd199, 32'd4341},
{32'd1429, 32'd2783, 32'd5847, 32'd161},
{-32'd3703, 32'd1293, -32'd7617, -32'd3107},
{-32'd844, -32'd4097, -32'd6569, 32'd1382},
{-32'd2922, 32'd1903, -32'd557, -32'd2125},
{32'd2639, -32'd7013, -32'd3357, -32'd673},
{32'd607, -32'd22, -32'd8826, -32'd4205},
{-32'd9011, -32'd3995, -32'd939, -32'd965},
{32'd40, 32'd584, 32'd799, 32'd4305},
{32'd3481, -32'd968, 32'd2204, -32'd904},
{-32'd3429, 32'd3529, -32'd1898, -32'd3675},
{32'd4786, 32'd9693, -32'd5989, 32'd1976},
{-32'd1480, -32'd5382, 32'd2498, 32'd2883},
{32'd11347, -32'd746, -32'd2466, 32'd3254},
{32'd676, -32'd3202, 32'd3662, -32'd99},
{-32'd11750, 32'd879, -32'd11940, -32'd3902},
{-32'd1088, 32'd1261, 32'd5254, 32'd1049},
{-32'd6917, -32'd5784, 32'd5468, -32'd6079},
{32'd10655, 32'd1565, 32'd3540, 32'd7993},
{-32'd4261, 32'd3210, -32'd4237, -32'd3382},
{32'd7348, 32'd997, -32'd1326, 32'd2958},
{32'd3276, 32'd1800, 32'd1132, -32'd3297},
{32'd7883, 32'd5685, -32'd2162, 32'd7554},
{-32'd1394, -32'd4480, 32'd11734, -32'd3285},
{32'd174, 32'd3031, 32'd3168, 32'd723},
{32'd6281, 32'd1257, -32'd2060, -32'd580},
{32'd5027, 32'd7411, 32'd1414, -32'd2684},
{-32'd6869, -32'd465, 32'd569, -32'd8035},
{-32'd3054, 32'd4168, -32'd1122, 32'd6254},
{-32'd1072, 32'd0, 32'd1519, -32'd4668},
{-32'd5785, -32'd4558, -32'd3642, 32'd1338},
{-32'd7288, -32'd3451, -32'd18, -32'd3818},
{32'd5216, 32'd3665, -32'd2511, 32'd15},
{-32'd178, -32'd1830, 32'd2486, -32'd3064},
{-32'd1651, 32'd676, -32'd789, -32'd655},
{-32'd2684, 32'd1277, 32'd1974, -32'd3453},
{32'd1223, -32'd2014, -32'd5157, -32'd161},
{32'd4047, 32'd5248, 32'd530, 32'd4653},
{32'd9221, 32'd5991, 32'd9657, -32'd2728},
{32'd2597, 32'd5679, 32'd2602, 32'd249},
{32'd2342, -32'd3608, 32'd3698, 32'd3910},
{-32'd4403, 32'd5019, -32'd4595, -32'd1657},
{-32'd6176, -32'd1586, 32'd9850, -32'd1039},
{32'd2602, -32'd2583, -32'd1861, 32'd2123},
{-32'd2026, -32'd1259, -32'd3261, -32'd4531},
{32'd930, -32'd4960, -32'd875, 32'd2685},
{-32'd2559, 32'd548, -32'd10085, -32'd7167},
{32'd4435, 32'd3062, -32'd3891, 32'd794},
{-32'd3259, 32'd2247, 32'd6717, -32'd927},
{32'd5590, 32'd4981, -32'd3533, 32'd3918},
{-32'd7411, -32'd1682, 32'd3353, -32'd3810},
{-32'd494, 32'd10685, -32'd1247, -32'd3030},
{-32'd2539, 32'd1302, 32'd1335, -32'd859},
{32'd1904, -32'd2835, -32'd5155, 32'd1627},
{32'd1418, 32'd427, 32'd4566, -32'd3839},
{32'd1502, 32'd6397, -32'd1983, -32'd984},
{-32'd2957, -32'd669, 32'd232, -32'd220},
{-32'd12163, 32'd4664, 32'd459, 32'd1153},
{-32'd634, -32'd1199, -32'd56, 32'd3687},
{-32'd827, 32'd4395, 32'd6330, -32'd2231},
{32'd1240, -32'd11880, -32'd1114, 32'd1835},
{-32'd3715, 32'd2721, 32'd3935, 32'd288},
{32'd3803, 32'd6188, -32'd2858, -32'd1861},
{32'd9457, -32'd1649, 32'd2421, 32'd1605},
{-32'd674, 32'd1122, 32'd2516, -32'd766},
{-32'd1417, 32'd8194, -32'd1023, 32'd3789},
{-32'd1403, -32'd5329, 32'd3209, 32'd4043},
{-32'd12508, 32'd68, -32'd227, -32'd5090},
{-32'd1040, 32'd4046, 32'd2881, 32'd2790},
{32'd9206, 32'd5347, -32'd1200, -32'd285},
{-32'd442, -32'd2807, -32'd9088, 32'd7802},
{-32'd4272, -32'd3150, -32'd2279, -32'd2909},
{-32'd9028, -32'd7894, 32'd811, 32'd1154},
{32'd2060, -32'd2031, 32'd3356, -32'd3857},
{32'd653, 32'd4583, 32'd2793, 32'd4580},
{-32'd4503, 32'd6338, -32'd6014, -32'd1773},
{32'd9927, 32'd6688, 32'd2778, 32'd3493},
{-32'd2133, 32'd6080, 32'd938, 32'd2260},
{32'd23, 32'd1658, -32'd2870, 32'd4398},
{32'd1687, -32'd6474, -32'd9912, 32'd1472},
{32'd5360, 32'd2640, 32'd3280, 32'd4203},
{-32'd1628, 32'd914, -32'd3918, 32'd1290},
{-32'd6827, -32'd1013, 32'd6362, 32'd454},
{32'd9324, 32'd2322, 32'd419, 32'd5301},
{-32'd5614, -32'd2420, 32'd588, -32'd4682},
{-32'd11918, -32'd3966, 32'd357, -32'd1310},
{-32'd7420, 32'd4564, 32'd4340, -32'd5680},
{-32'd1803, 32'd4408, -32'd3543, -32'd1163},
{32'd1717, -32'd6393, -32'd5389, 32'd4887},
{-32'd1180, 32'd4221, 32'd1836, 32'd858},
{-32'd3562, -32'd1346, 32'd4810, -32'd7983},
{32'd4111, -32'd5845, 32'd2640, -32'd971},
{32'd6206, 32'd1538, 32'd12056, -32'd1045},
{-32'd5173, -32'd3977, -32'd3080, -32'd724},
{-32'd4431, 32'd9494, 32'd4441, 32'd4789},
{32'd510, -32'd5488, 32'd13, 32'd1838},
{32'd5959, 32'd3305, -32'd3476, 32'd2352},
{-32'd2848, 32'd4518, 32'd2315, 32'd2671},
{-32'd5561, 32'd358, -32'd5424, 32'd787},
{32'd253, -32'd4784, -32'd12932, -32'd5747},
{-32'd4672, 32'd5464, 32'd7989, 32'd4197},
{-32'd4667, 32'd3437, -32'd1034, -32'd7134},
{-32'd7667, 32'd10483, -32'd1081, -32'd6034},
{32'd874, 32'd9947, -32'd3199, 32'd8295},
{32'd12728, 32'd3275, -32'd1458, 32'd1271},
{-32'd9809, -32'd1158, -32'd522, 32'd1896},
{-32'd3584, 32'd4242, -32'd2748, -32'd6281},
{32'd2572, -32'd11698, -32'd10018, 32'd1407},
{32'd1256, -32'd5833, 32'd3534, 32'd7088},
{32'd5333, 32'd3582, -32'd2, 32'd3183},
{-32'd180, 32'd2152, 32'd6851, 32'd2764},
{32'd252, 32'd238, -32'd5465, 32'd724},
{-32'd1414, -32'd5694, 32'd4756, 32'd878},
{32'd1263, 32'd4243, 32'd1703, 32'd2857},
{-32'd4523, -32'd8, -32'd729, -32'd1953},
{-32'd7437, -32'd5351, 32'd4609, -32'd4072},
{-32'd8254, -32'd2991, -32'd3987, -32'd3063},
{-32'd2279, -32'd4745, 32'd1198, 32'd1275},
{32'd1150, 32'd5892, -32'd3134, -32'd7111},
{-32'd1413, -32'd2813, -32'd5125, 32'd1569},
{32'd7351, -32'd1528, -32'd6796, -32'd3513},
{-32'd4500, 32'd918, -32'd190, -32'd1517},
{-32'd296, 32'd1535, -32'd1511, 32'd6022},
{32'd391, -32'd8777, -32'd690, 32'd146},
{-32'd835, 32'd412, -32'd4509, 32'd1083},
{32'd1294, -32'd5337, -32'd370, -32'd3193},
{-32'd177, 32'd10881, -32'd8766, -32'd1352},
{-32'd5510, 32'd4346, -32'd383, -32'd1401},
{32'd6722, -32'd2721, -32'd691, 32'd6237},
{32'd1288, 32'd2107, -32'd6046, 32'd1077},
{-32'd1885, -32'd6479, 32'd5234, -32'd3541},
{-32'd1629, 32'd7371, 32'd2038, -32'd368},
{32'd5894, -32'd3249, -32'd1708, 32'd2681},
{32'd3428, -32'd1060, -32'd719, 32'd3725},
{-32'd11949, -32'd3432, 32'd3043, -32'd7074},
{-32'd3878, -32'd617, -32'd1688, -32'd5677},
{-32'd655, -32'd1086, 32'd3709, -32'd485},
{32'd13005, -32'd6323, 32'd422, 32'd1494},
{-32'd5631, -32'd1729, 32'd1989, -32'd7993},
{-32'd1431, 32'd4198, -32'd1586, 32'd1623},
{32'd4900, 32'd18, -32'd5910, -32'd1814},
{-32'd1348, 32'd3565, -32'd3781, 32'd4808},
{-32'd1956, 32'd600, 32'd4384, 32'd1696},
{32'd5016, 32'd2294, -32'd470, 32'd2743},
{-32'd5099, 32'd3804, -32'd13028, -32'd973},
{32'd4023, 32'd1401, 32'd4482, -32'd408},
{32'd845, -32'd2619, -32'd2774, 32'd169},
{-32'd6056, 32'd737, 32'd6188, -32'd1861},
{-32'd1987, -32'd1642, -32'd3097, 32'd3811},
{-32'd5978, -32'd2497, -32'd458, -32'd4433},
{-32'd5362, -32'd2894, 32'd3724, -32'd7569},
{32'd4545, 32'd2601, -32'd6372, -32'd168},
{-32'd1306, -32'd5982, 32'd4546, -32'd8070},
{-32'd4560, -32'd1926, 32'd1495, -32'd663},
{32'd135, -32'd4363, 32'd3076, 32'd289},
{-32'd3130, -32'd2903, 32'd225, 32'd1998},
{32'd7589, 32'd4090, 32'd1307, 32'd3322},
{-32'd5414, -32'd1856, 32'd269, 32'd837},
{32'd1932, 32'd3731, -32'd2796, 32'd855},
{-32'd5307, -32'd5716, 32'd7936, 32'd1689},
{-32'd2187, -32'd5266, 32'd8938, 32'd1456},
{32'd3996, -32'd4065, -32'd2676, -32'd2014},
{-32'd6976, 32'd2732, -32'd6975, 32'd5777},
{-32'd4478, 32'd7049, -32'd3459, -32'd2262},
{-32'd2815, 32'd677, -32'd2892, -32'd6537},
{-32'd1575, 32'd5093, 32'd5123, -32'd3482},
{-32'd1211, -32'd647, 32'd1092, -32'd7714},
{-32'd2891, 32'd1261, 32'd8309, -32'd3434},
{-32'd6915, -32'd2899, 32'd4018, 32'd2603},
{32'd5438, 32'd16108, 32'd1530, -32'd2185},
{32'd4115, 32'd2995, -32'd308, -32'd3575},
{32'd758, 32'd6185, 32'd6789, 32'd2761},
{32'd3804, -32'd9311, -32'd3073, -32'd5942},
{-32'd483, -32'd3826, -32'd601, -32'd2435},
{-32'd7854, -32'd4115, -32'd1111, -32'd6152},
{32'd2732, -32'd2389, -32'd3498, -32'd7718},
{-32'd1654, 32'd267, 32'd1685, -32'd680},
{32'd7260, -32'd3819, -32'd10510, 32'd2617},
{32'd3308, 32'd721, 32'd5929, 32'd5530},
{32'd3485, 32'd7798, -32'd1630, 32'd4990},
{-32'd7185, 32'd10353, 32'd6746, -32'd1464},
{32'd10874, -32'd48, 32'd10246, 32'd580},
{32'd3128, -32'd678, -32'd3467, 32'd3687},
{-32'd6292, 32'd3652, -32'd2819, -32'd830},
{-32'd11300, -32'd6268, -32'd1323, -32'd6404},
{32'd3582, 32'd47, 32'd3798, -32'd559},
{-32'd3673, -32'd1016, -32'd11181, -32'd30},
{-32'd287, -32'd1431, -32'd4660, -32'd3351},
{-32'd1102, -32'd8708, -32'd2185, 32'd2052},
{32'd4155, 32'd8011, -32'd1455, 32'd4960},
{32'd6370, 32'd2296, 32'd5298, 32'd4269},
{32'd1078, 32'd4087, -32'd6943, 32'd3064},
{32'd2932, -32'd6048, 32'd7421, 32'd1399},
{32'd1658, -32'd6527, -32'd577, -32'd758},
{32'd1779, 32'd1094, 32'd3775, 32'd2188},
{32'd6261, 32'd90, -32'd3609, 32'd5381},
{32'd884, 32'd7022, -32'd69, -32'd3637},
{32'd1581, 32'd3594, 32'd1702, -32'd165},
{32'd1595, -32'd2916, 32'd4960, -32'd7187},
{-32'd6957, -32'd1491, -32'd8050, -32'd6190},
{32'd1473, 32'd764, -32'd4136, -32'd4661},
{-32'd697, 32'd158, -32'd1830, 32'd118},
{-32'd1567, -32'd11591, 32'd4786, -32'd411},
{32'd3246, 32'd4320, -32'd4840, -32'd2004},
{-32'd2219, 32'd951, -32'd2811, -32'd2519},
{-32'd2156, -32'd451, -32'd3767, -32'd3708},
{-32'd580, -32'd269, 32'd2707, 32'd3733},
{32'd382, -32'd151, 32'd6945, -32'd3286},
{-32'd3363, -32'd10108, 32'd7947, -32'd913},
{-32'd9655, -32'd1651, -32'd749, 32'd4352},
{-32'd1243, 32'd2837, 32'd580, -32'd6424},
{-32'd445, 32'd6595, -32'd5118, -32'd360},
{-32'd4826, -32'd2248, 32'd2216, -32'd3215},
{32'd8457, 32'd4823, -32'd4538, -32'd52},
{32'd500, -32'd9340, 32'd4280, -32'd2197},
{-32'd7803, 32'd10151, 32'd2325, -32'd2106},
{32'd1053, 32'd10612, -32'd567, -32'd2124},
{32'd1957, 32'd2895, -32'd2220, 32'd2722},
{32'd1065, -32'd1171, -32'd2686, -32'd7474},
{32'd7460, 32'd5012, -32'd2408, -32'd1940},
{-32'd3609, -32'd2206, -32'd1289, 32'd2166},
{-32'd6100, -32'd128, 32'd1577, -32'd2592},
{-32'd219, -32'd49, 32'd3092, -32'd4612},
{32'd2679, -32'd328, -32'd8404, -32'd699},
{32'd2496, -32'd104, -32'd5392, 32'd2936},
{32'd6279, -32'd3467, -32'd2095, 32'd4351},
{-32'd5526, 32'd1172, 32'd2542, -32'd5833},
{-32'd1030, -32'd2813, 32'd1532, 32'd1308},
{32'd7280, 32'd5985, 32'd4353, 32'd8589},
{-32'd923, -32'd5620, -32'd2362, 32'd3302},
{32'd3104, -32'd6057, 32'd1029, -32'd454},
{32'd6979, -32'd4849, -32'd1867, 32'd5204},
{-32'd3903, -32'd4450, 32'd5246, 32'd1056},
{32'd5615, -32'd5002, 32'd674, 32'd2412},
{32'd608, -32'd604, 32'd6298, 32'd330},
{-32'd1873, 32'd1054, -32'd5357, 32'd1917},
{32'd2570, -32'd3295, -32'd4380, 32'd742},
{32'd5686, 32'd687, -32'd220, -32'd2472},
{-32'd381, 32'd1711, -32'd6512, -32'd7493},
{-32'd4545, -32'd6420, -32'd8508, -32'd4424},
{32'd7659, 32'd6317, 32'd5154, 32'd3541},
{32'd2379, 32'd642, 32'd6945, 32'd4174},
{-32'd4802, -32'd4579, -32'd822, -32'd2064},
{-32'd803, 32'd4285, -32'd1819, 32'd1160},
{32'd2898, 32'd6963, -32'd3815, 32'd6650},
{-32'd3237, 32'd775, 32'd4842, 32'd6158},
{-32'd3583, -32'd5505, -32'd5455, 32'd297},
{32'd4129, -32'd6423, 32'd3927, 32'd5871},
{-32'd3123, 32'd4336, -32'd5148, -32'd211},
{-32'd1249, 32'd5150, -32'd1396, 32'd2691},
{-32'd6051, 32'd4729, 32'd3672, 32'd68},
{32'd6520, 32'd4664, -32'd6804, 32'd161},
{32'd3203, -32'd5318, -32'd9501, 32'd580},
{32'd2429, -32'd4435, -32'd6163, 32'd3479},
{32'd209, 32'd3212, 32'd24, -32'd804},
{32'd833, 32'd6991, 32'd1569, 32'd4836},
{-32'd2925, 32'd5786, 32'd4283, -32'd5823},
{32'd2116, 32'd1702, -32'd470, -32'd5098},
{-32'd734, 32'd8303, 32'd1703, 32'd4374},
{-32'd631, -32'd3344, 32'd3219, -32'd3473},
{32'd12287, 32'd6094, 32'd993, 32'd6929},
{32'd401, -32'd4714, 32'd5023, -32'd81},
{-32'd6510, 32'd1656, -32'd753, -32'd4582},
{32'd1977, -32'd5023, 32'd865, -32'd6060},
{32'd10576, 32'd4227, -32'd3651, 32'd3500},
{32'd3246, 32'd1927, -32'd6634, 32'd1129},
{32'd3149, 32'd6587, 32'd1672, 32'd1485},
{32'd5221, -32'd446, -32'd3263, -32'd7178},
{32'd2081, 32'd3532, -32'd2232, 32'd6048},
{-32'd4527, -32'd8046, -32'd4870, -32'd1340},
{32'd3723, 32'd7871, -32'd5252, 32'd4709},
{-32'd900, 32'd520, 32'd580, -32'd1536},
{-32'd5659, -32'd3904, -32'd13469, -32'd3800},
{-32'd3985, 32'd1723, -32'd8418, 32'd5408},
{-32'd6742, 32'd814, 32'd2275, 32'd2019},
{32'd1065, 32'd5693, 32'd1320, 32'd5228},
{32'd6329, -32'd655, 32'd7006, 32'd973},
{-32'd4403, -32'd2143, -32'd4752, 32'd1096},
{32'd2058, -32'd10356, -32'd913, -32'd1947},
{-32'd3327, -32'd11948, 32'd5274, -32'd5377},
{-32'd9467, 32'd425, -32'd5295, -32'd3474},
{32'd5625, 32'd1767, -32'd7369, 32'd3270},
{32'd241, -32'd1771, -32'd5027, 32'd2659},
{-32'd5399, 32'd2398, -32'd5703, -32'd3572}
},
{{-32'd5637, 32'd3997, 32'd10484, 32'd2891},
{-32'd6479, -32'd13429, 32'd2427, 32'd10636},
{-32'd8690, 32'd2912, 32'd2045, -32'd3613},
{-32'd4312, -32'd5586, 32'd1378, 32'd4025},
{-32'd13712, 32'd5977, 32'd7663, 32'd6064},
{32'd5958, -32'd6378, 32'd4580, 32'd4267},
{32'd5250, 32'd7331, -32'd7701, 32'd7366},
{32'd4000, -32'd3042, 32'd749, -32'd6928},
{32'd114, 32'd1428, 32'd11000, -32'd9444},
{32'd2322, 32'd4966, 32'd5630, -32'd979},
{-32'd11707, -32'd663, -32'd4095, -32'd951},
{32'd1827, -32'd6040, -32'd1462, -32'd947},
{32'd7822, 32'd13310, -32'd1523, 32'd4263},
{32'd14107, -32'd4209, -32'd5184, -32'd5236},
{32'd13400, -32'd13729, -32'd8270, -32'd17142},
{32'd15751, -32'd1708, 32'd5367, 32'd1376},
{32'd3010, 32'd7556, 32'd648, 32'd3486},
{32'd15732, -32'd828, -32'd7653, -32'd8983},
{-32'd18879, -32'd2979, 32'd4093, -32'd4190},
{-32'd13820, 32'd19495, -32'd2976, -32'd3634},
{-32'd5125, -32'd2447, 32'd7091, 32'd13197},
{32'd957, -32'd1062, -32'd5595, -32'd10383},
{-32'd5323, -32'd1060, -32'd212, 32'd441},
{32'd677, -32'd12454, -32'd6037, -32'd2362},
{-32'd2139, -32'd4547, -32'd1273, 32'd263},
{32'd2924, -32'd7292, 32'd3204, -32'd1026},
{-32'd13187, 32'd375, 32'd3594, -32'd12257},
{32'd540, 32'd2445, 32'd7143, -32'd2772},
{32'd21679, -32'd6462, 32'd10791, -32'd2663},
{-32'd1927, 32'd6011, -32'd10876, -32'd3261},
{32'd290, -32'd13955, 32'd973, 32'd4721},
{32'd5418, -32'd8997, -32'd744, -32'd13582},
{32'd3649, 32'd6320, 32'd3558, -32'd1471},
{32'd527, -32'd5871, 32'd5673, -32'd4989},
{32'd3546, 32'd5979, -32'd1966, 32'd2792},
{-32'd5374, -32'd19249, 32'd5610, 32'd7841},
{32'd7675, 32'd4337, -32'd900, -32'd9056},
{32'd10934, -32'd4544, 32'd8699, 32'd7383},
{32'd2798, -32'd1661, 32'd5713, -32'd780},
{-32'd5832, -32'd3321, -32'd8536, 32'd3146},
{32'd8289, -32'd9952, 32'd5974, 32'd19472},
{-32'd2333, -32'd5949, -32'd2850, 32'd7216},
{32'd11832, -32'd996, -32'd4876, 32'd4801},
{32'd6541, -32'd6668, -32'd9157, 32'd677},
{32'd8619, 32'd959, -32'd9420, -32'd19826},
{-32'd7019, 32'd2326, -32'd302, 32'd5040},
{-32'd2842, 32'd5957, -32'd15365, -32'd2932},
{32'd2142, -32'd6576, -32'd8544, -32'd10574},
{-32'd1674, 32'd6690, -32'd4407, -32'd7448},
{-32'd4676, -32'd211, 32'd7364, -32'd162},
{-32'd3578, 32'd13597, -32'd3686, -32'd13069},
{32'd6334, -32'd25, -32'd6752, -32'd4479},
{-32'd16339, -32'd8763, 32'd323, 32'd1516},
{-32'd7473, 32'd6648, 32'd657, 32'd6317},
{32'd10977, 32'd367, 32'd10442, 32'd2922},
{-32'd2658, -32'd3931, -32'd6461, -32'd504},
{-32'd8801, 32'd7235, -32'd1419, 32'd9456},
{32'd8230, -32'd3642, -32'd14703, -32'd6531},
{32'd1717, -32'd5316, -32'd4345, -32'd680},
{-32'd12528, -32'd10091, 32'd31, 32'd3964},
{-32'd10282, -32'd1377, 32'd11652, 32'd2875},
{-32'd4072, 32'd7029, 32'd3307, 32'd8642},
{32'd528, -32'd4478, -32'd2814, -32'd10625},
{-32'd9185, 32'd1060, -32'd2128, 32'd4376},
{-32'd2687, 32'd637, 32'd361, -32'd4792},
{-32'd6805, -32'd271, 32'd871, -32'd465},
{32'd3437, -32'd9349, 32'd5785, 32'd8640},
{-32'd6854, -32'd5309, 32'd3679, -32'd2810},
{-32'd631, -32'd3318, 32'd2032, -32'd5510},
{-32'd5153, 32'd1019, -32'd6984, -32'd8153},
{32'd3314, -32'd3546, 32'd2835, -32'd3008},
{32'd177, -32'd7826, -32'd1251, -32'd4024},
{32'd5365, 32'd101, -32'd415, 32'd1111},
{-32'd17832, -32'd141, 32'd2411, 32'd2977},
{32'd5074, 32'd5714, 32'd13453, 32'd1648},
{32'd22063, -32'd3772, -32'd9032, 32'd14742},
{32'd8231, 32'd9152, -32'd5379, 32'd1008},
{32'd5108, -32'd11446, -32'd2510, -32'd1229},
{-32'd825, 32'd3992, 32'd3266, 32'd5588},
{-32'd1618, -32'd15506, -32'd13433, -32'd2217},
{-32'd3775, 32'd7964, 32'd2223, -32'd6038},
{-32'd11981, 32'd6249, -32'd6204, 32'd6380},
{-32'd1728, -32'd275, 32'd4233, 32'd6942},
{32'd12326, 32'd11328, 32'd14920, 32'd5648},
{-32'd3862, -32'd3718, -32'd1453, -32'd9702},
{-32'd1126, -32'd9598, -32'd5531, 32'd1340},
{32'd282, 32'd14245, 32'd1284, 32'd3483},
{-32'd2898, -32'd8252, -32'd50, -32'd624},
{-32'd2521, 32'd5250, -32'd4266, -32'd3307},
{32'd3127, -32'd8214, 32'd5100, -32'd10113},
{32'd3973, -32'd1384, 32'd8176, 32'd5340},
{-32'd12758, 32'd5553, -32'd141, 32'd6074},
{-32'd12570, -32'd2078, -32'd14365, -32'd18737},
{32'd6979, 32'd8591, 32'd109, 32'd9674},
{32'd16542, 32'd2188, -32'd7093, 32'd3118},
{32'd4580, 32'd8607, -32'd7693, 32'd5656},
{32'd1468, 32'd3116, 32'd3016, -32'd6551},
{32'd8534, -32'd8367, 32'd4842, -32'd3232},
{32'd4263, 32'd4023, 32'd4378, 32'd6836},
{32'd9292, 32'd9907, 32'd10131, -32'd4150},
{32'd3035, -32'd10115, 32'd120, 32'd8865},
{32'd1944, -32'd8019, -32'd6463, 32'd2781},
{-32'd75, 32'd7334, 32'd1672, 32'd2689},
{-32'd3628, 32'd3943, 32'd5875, 32'd3157},
{-32'd1562, -32'd2736, -32'd4044, -32'd2837},
{-32'd5303, 32'd3331, 32'd2908, 32'd70},
{32'd15990, 32'd7228, -32'd2664, -32'd321},
{32'd1535, -32'd11, 32'd8285, -32'd3234},
{-32'd5436, 32'd597, 32'd7416, -32'd4218},
{-32'd6300, -32'd4407, 32'd3226, -32'd53},
{-32'd10483, 32'd1737, -32'd8985, -32'd13784},
{32'd3581, 32'd3514, -32'd966, 32'd1385},
{-32'd6613, 32'd7629, 32'd2760, 32'd3457},
{32'd2009, 32'd9738, -32'd533, -32'd9567},
{32'd2850, 32'd5340, 32'd7836, 32'd4684},
{-32'd1647, -32'd4249, 32'd4968, -32'd584},
{32'd3896, 32'd2388, 32'd7467, 32'd506},
{32'd5390, -32'd7207, -32'd3899, -32'd12432},
{32'd10817, 32'd2951, -32'd1826, -32'd13949},
{32'd2361, -32'd218, 32'd554, 32'd3349},
{-32'd15242, 32'd3621, 32'd4041, 32'd7657},
{-32'd6334, 32'd1426, -32'd6535, -32'd8361},
{-32'd6882, -32'd9415, -32'd5696, 32'd3567},
{32'd9182, -32'd5996, -32'd1049, -32'd1994},
{-32'd14469, 32'd1115, -32'd792, 32'd510},
{32'd9057, 32'd14592, 32'd5378, -32'd1561},
{32'd2911, -32'd19137, -32'd1875, -32'd2315},
{32'd3924, -32'd15550, 32'd1680, 32'd1962},
{32'd6412, 32'd5765, -32'd315, -32'd6248},
{-32'd6187, -32'd2858, 32'd11132, -32'd1116},
{-32'd12678, -32'd373, -32'd5262, -32'd3632},
{-32'd8725, -32'd4458, -32'd8260, -32'd7717},
{-32'd8000, -32'd1868, -32'd15549, -32'd1761},
{32'd4749, 32'd634, 32'd5584, -32'd2312},
{-32'd8760, -32'd5712, 32'd12125, -32'd868},
{32'd5667, -32'd1047, -32'd8532, -32'd10891},
{-32'd6078, 32'd7432, 32'd3387, -32'd8392},
{-32'd6565, -32'd8005, 32'd439, 32'd8922},
{32'd6095, -32'd4541, -32'd1331, 32'd2888},
{32'd5197, -32'd4629, -32'd289, 32'd874},
{-32'd8595, -32'd3324, 32'd7596, 32'd2463},
{32'd788, 32'd7459, -32'd7126, 32'd221},
{32'd8035, -32'd11220, 32'd4005, 32'd12216},
{32'd4319, 32'd12558, 32'd3600, 32'd1060},
{-32'd3823, -32'd3457, -32'd2556, -32'd2443},
{32'd6809, 32'd3497, -32'd436, -32'd1788},
{-32'd11776, 32'd4887, -32'd6421, 32'd5904},
{-32'd10516, 32'd1120, -32'd5327, 32'd5711},
{32'd3164, -32'd8655, -32'd5854, 32'd5083},
{-32'd8740, -32'd16020, -32'd16320, -32'd5330},
{32'd2915, 32'd6818, -32'd205, -32'd3403},
{-32'd5142, 32'd15582, 32'd4450, 32'd9540},
{-32'd2744, 32'd654, 32'd8356, 32'd9429},
{32'd11319, 32'd12156, -32'd9694, 32'd5909},
{-32'd14728, 32'd1088, -32'd4536, -32'd11005},
{-32'd2994, -32'd3632, 32'd3765, -32'd4201},
{-32'd9246, 32'd5709, 32'd2532, 32'd5522},
{32'd4014, -32'd2020, -32'd1878, 32'd2326},
{32'd7411, 32'd5101, 32'd7706, 32'd3856},
{32'd5286, 32'd8987, 32'd11031, -32'd5078},
{-32'd10361, -32'd4400, 32'd5098, -32'd18982},
{32'd226, -32'd3502, 32'd7495, -32'd5812},
{-32'd9782, 32'd4648, -32'd6013, -32'd3786},
{32'd7098, 32'd5985, 32'd4623, 32'd11428},
{32'd8574, -32'd1331, 32'd14738, 32'd13257},
{-32'd8665, -32'd4652, -32'd3249, 32'd1510},
{-32'd1633, 32'd4158, 32'd3406, -32'd4804},
{32'd4806, -32'd5295, -32'd16949, -32'd3550},
{32'd12376, 32'd4073, 32'd3951, 32'd3138},
{-32'd3269, -32'd5474, -32'd4123, -32'd4898},
{32'd4656, -32'd12402, 32'd925, -32'd9676},
{-32'd13916, 32'd1586, -32'd8639, -32'd6001},
{32'd4350, 32'd1038, 32'd2582, 32'd4350},
{-32'd10733, 32'd2764, -32'd6354, -32'd12737},
{32'd3075, -32'd2203, 32'd144, -32'd4922},
{-32'd4947, -32'd3908, -32'd1100, -32'd8111},
{32'd8614, -32'd2184, -32'd4899, 32'd9578},
{-32'd962, 32'd1981, 32'd7239, 32'd8863},
{32'd8021, -32'd1056, 32'd4752, -32'd2270},
{32'd724, 32'd5359, -32'd5941, -32'd12048},
{-32'd905, -32'd10856, 32'd4589, -32'd4368},
{32'd2503, 32'd1645, -32'd6142, -32'd33},
{32'd1569, -32'd20355, 32'd8001, 32'd10399},
{-32'd5165, 32'd13134, -32'd245, -32'd13005},
{32'd510, 32'd4311, -32'd183, -32'd7707},
{-32'd7542, 32'd4691, 32'd4881, 32'd5956},
{32'd7125, -32'd3669, 32'd975, -32'd2513},
{32'd2742, 32'd6782, 32'd6005, 32'd1017},
{32'd2927, 32'd7536, -32'd5468, 32'd2499},
{32'd4149, 32'd8675, 32'd4624, -32'd3796},
{32'd4198, -32'd2200, 32'd6704, 32'd603},
{-32'd3866, -32'd13795, -32'd2355, -32'd7402},
{32'd8739, -32'd5684, 32'd1562, -32'd4035},
{-32'd2673, -32'd7892, 32'd5367, -32'd2486},
{-32'd2358, -32'd7432, 32'd5221, -32'd4089},
{-32'd14739, -32'd7000, -32'd9374, -32'd2079},
{-32'd15571, -32'd7519, -32'd2340, 32'd5929},
{-32'd8184, -32'd2379, 32'd9733, 32'd14961},
{-32'd1691, -32'd2071, -32'd398, -32'd5698},
{-32'd952, 32'd6639, 32'd12153, -32'd2765},
{-32'd7864, -32'd595, -32'd4710, -32'd9900},
{-32'd1258, -32'd6288, -32'd12460, -32'd8843},
{-32'd7534, 32'd8022, 32'd510, -32'd3070},
{32'd8615, 32'd3108, 32'd415, 32'd3365},
{-32'd1299, 32'd10454, 32'd7489, -32'd12337},
{32'd6466, -32'd5905, -32'd5374, 32'd9013},
{32'd7422, 32'd6968, 32'd409, 32'd9145},
{-32'd494, 32'd5171, 32'd3316, -32'd10904},
{32'd9341, 32'd11205, -32'd5636, -32'd3901},
{-32'd726, 32'd4550, 32'd8379, -32'd2368},
{32'd11196, -32'd5854, -32'd4243, 32'd9359},
{-32'd4965, 32'd4157, 32'd6417, -32'd2059},
{-32'd10199, 32'd226, 32'd4487, -32'd7464},
{-32'd1643, -32'd11082, 32'd3970, 32'd745},
{-32'd8607, 32'd10739, -32'd2292, -32'd579},
{-32'd496, 32'd7079, 32'd55, -32'd9960},
{-32'd1960, 32'd9265, 32'd11309, -32'd12483},
{32'd7661, 32'd1478, -32'd8959, -32'd6548},
{32'd8366, 32'd10189, 32'd9848, 32'd15052},
{32'd12945, 32'd1636, -32'd2481, -32'd5034},
{32'd3501, 32'd9611, -32'd411, 32'd664},
{-32'd7410, 32'd391, -32'd1641, -32'd7195},
{32'd5323, 32'd4556, 32'd3632, 32'd480},
{32'd6469, 32'd5528, -32'd3059, -32'd4791},
{32'd2286, 32'd1340, 32'd1314, 32'd12489},
{32'd5308, -32'd5997, 32'd9937, 32'd3548},
{-32'd3435, -32'd4307, 32'd7707, -32'd10261},
{-32'd4636, -32'd13713, 32'd10854, 32'd1726},
{32'd11478, 32'd10085, -32'd4017, 32'd902},
{32'd3144, 32'd4862, 32'd4742, -32'd20908},
{-32'd1752, -32'd7119, -32'd948, 32'd214},
{-32'd8721, 32'd2456, -32'd128, -32'd3157},
{-32'd2521, -32'd7639, 32'd3868, 32'd6600},
{-32'd4755, -32'd376, -32'd357, -32'd416},
{32'd14967, 32'd7288, -32'd2278, -32'd10237},
{-32'd897, -32'd1061, -32'd3009, -32'd6757},
{-32'd6317, 32'd6751, 32'd882, 32'd12732},
{32'd10397, 32'd4529, -32'd7609, 32'd2955},
{-32'd7548, -32'd7546, 32'd16116, 32'd13167},
{32'd8016, -32'd3229, -32'd1650, 32'd3833},
{-32'd3452, -32'd6424, -32'd1847, 32'd9370},
{32'd6660, -32'd718, 32'd739, 32'd1567},
{-32'd2047, -32'd9247, 32'd237, 32'd3103},
{32'd7221, 32'd12024, 32'd6189, 32'd1582},
{32'd9616, 32'd11824, 32'd7393, 32'd896},
{-32'd11173, -32'd2528, -32'd10166, -32'd1768},
{32'd12108, 32'd10375, -32'd4599, -32'd5760},
{-32'd11225, -32'd2672, -32'd3896, -32'd10183},
{32'd17120, 32'd568, -32'd1016, 32'd7222},
{32'd9390, 32'd6389, 32'd13673, 32'd10688},
{-32'd7878, -32'd4848, 32'd1748, 32'd7903},
{32'd2653, -32'd8053, -32'd7997, -32'd3542},
{-32'd1557, 32'd7539, 32'd450, -32'd2606},
{-32'd3782, 32'd7549, -32'd10699, -32'd1398},
{32'd1050, 32'd10333, -32'd7935, -32'd2973},
{32'd9375, 32'd5554, 32'd2305, 32'd198},
{-32'd10629, 32'd16388, -32'd3654, 32'd4640},
{32'd2800, 32'd7923, 32'd6398, 32'd2669},
{32'd7746, -32'd1790, -32'd11239, -32'd8126},
{32'd11702, 32'd8626, 32'd9355, -32'd2253},
{32'd11264, -32'd5569, -32'd4782, -32'd7234},
{32'd22036, -32'd7055, 32'd7906, 32'd5019},
{-32'd6445, -32'd4780, -32'd7778, 32'd11597},
{32'd7998, 32'd4583, -32'd10841, -32'd11709},
{-32'd4479, 32'd42, 32'd3095, -32'd13247},
{32'd10143, -32'd8499, -32'd2174, -32'd72},
{32'd18612, 32'd5458, 32'd2194, -32'd4320},
{-32'd744, -32'd1947, -32'd3364, 32'd1585},
{32'd6502, -32'd12441, -32'd2516, -32'd11003},
{-32'd324, -32'd3646, -32'd2083, 32'd760},
{-32'd4137, -32'd7596, 32'd3586, 32'd1575},
{-32'd15762, 32'd392, -32'd3113, -32'd3692},
{-32'd2899, -32'd2951, -32'd6201, 32'd3337},
{-32'd4612, 32'd197, -32'd5258, -32'd514},
{-32'd3441, 32'd1064, -32'd3646, -32'd6983},
{-32'd1319, -32'd2712, 32'd2855, -32'd796},
{32'd2173, 32'd4719, 32'd8394, -32'd60},
{32'd2825, -32'd6230, 32'd3110, 32'd6733},
{32'd3805, -32'd9307, 32'd1286, 32'd2453},
{-32'd7152, -32'd4861, -32'd1756, 32'd801},
{-32'd6450, -32'd7507, 32'd8718, -32'd7406},
{32'd5629, 32'd13462, -32'd10396, 32'd3583},
{32'd14481, -32'd97, 32'd4663, 32'd3376},
{-32'd3787, -32'd1715, -32'd4761, -32'd3462},
{32'd4866, -32'd10185, 32'd15275, 32'd13680},
{-32'd1691, 32'd3987, 32'd956, 32'd1190},
{-32'd7320, 32'd4324, -32'd1979, 32'd3117},
{-32'd1692, 32'd8979, -32'd3767, -32'd14600},
{-32'd85, 32'd9535, 32'd10833, 32'd4630},
{-32'd4011, -32'd9563, -32'd4020, -32'd2016},
{32'd291, 32'd5569, -32'd2232, 32'd5656},
{32'd2884, 32'd2924, -32'd5050, 32'd5781},
{32'd9187, 32'd182, 32'd16177, 32'd4416},
{32'd248, -32'd5612, 32'd3384, -32'd496},
{32'd649, -32'd1439, -32'd7924, -32'd121},
{32'd9131, 32'd10546, 32'd2915, -32'd2554},
{32'd2107, 32'd165, -32'd2366, -32'd136},
{32'd3646, -32'd4372, 32'd4409, -32'd717},
{-32'd9247, -32'd4350, 32'd2620, -32'd2908},
{-32'd1132, -32'd3745, 32'd8829, 32'd2082}
},
{{32'd5489, 32'd2836, -32'd195, 32'd5084},
{-32'd9013, -32'd7926, 32'd6048, -32'd13089},
{-32'd12645, 32'd2846, 32'd4564, -32'd4683},
{32'd3207, -32'd2134, 32'd1820, -32'd3493},
{-32'd9450, -32'd3664, -32'd5667, -32'd4154},
{32'd6503, -32'd6654, 32'd3090, -32'd385},
{32'd9105, 32'd938, 32'd12201, 32'd8630},
{32'd557, -32'd4749, 32'd3652, -32'd2218},
{32'd5309, 32'd621, 32'd10319, -32'd4733},
{32'd4338, 32'd13216, 32'd7353, 32'd214},
{-32'd9447, 32'd769, 32'd518, 32'd8610},
{32'd430, 32'd4747, 32'd3456, -32'd2297},
{-32'd675, -32'd799, -32'd8967, 32'd16147},
{32'd1115, 32'd246, -32'd6759, -32'd4780},
{-32'd9823, -32'd3306, -32'd4176, 32'd8754},
{32'd9305, 32'd1723, -32'd17981, 32'd116},
{32'd19139, 32'd127, -32'd954, 32'd11672},
{-32'd1478, 32'd2092, -32'd5674, 32'd6682},
{32'd268, -32'd8925, 32'd2849, -32'd1221},
{32'd8546, -32'd7318, 32'd9628, -32'd4396},
{-32'd24146, 32'd2709, 32'd7098, -32'd416},
{-32'd11846, -32'd8351, 32'd7379, 32'd2842},
{32'd10141, -32'd2227, -32'd1884, -32'd6381},
{-32'd10147, -32'd8579, -32'd5997, 32'd5293},
{32'd10865, 32'd4480, 32'd6123, 32'd10322},
{-32'd5383, -32'd5459, 32'd10870, -32'd1123},
{-32'd7458, -32'd3837, 32'd1027, -32'd4891},
{-32'd607, 32'd2584, 32'd3414, 32'd2480},
{-32'd1881, 32'd5354, 32'd1293, -32'd523},
{32'd2258, 32'd1043, 32'd1801, -32'd4076},
{32'd5694, -32'd6260, -32'd1517, -32'd319},
{32'd4061, -32'd7374, -32'd8715, -32'd19},
{32'd3948, -32'd687, -32'd2022, -32'd2415},
{-32'd11777, 32'd1317, -32'd7853, 32'd5743},
{32'd10202, 32'd7488, 32'd3217, 32'd925},
{32'd949, 32'd3253, 32'd11865, 32'd742},
{-32'd14088, -32'd8765, -32'd13650, 32'd95},
{32'd5599, 32'd2874, 32'd8361, -32'd521},
{-32'd1646, -32'd2594, 32'd5475, 32'd1312},
{32'd1459, 32'd17, -32'd3495, 32'd1738},
{-32'd13786, 32'd8874, -32'd5537, -32'd7889},
{32'd5027, 32'd7572, 32'd9265, 32'd6518},
{32'd19981, 32'd3057, -32'd766, 32'd13487},
{32'd5439, -32'd2166, -32'd6311, 32'd3266},
{-32'd3142, -32'd12232, -32'd5286, -32'd7286},
{-32'd2576, 32'd6993, 32'd4223, -32'd1699},
{32'd1170, -32'd7959, 32'd3638, 32'd6973},
{-32'd9210, -32'd8415, -32'd18286, 32'd3796},
{-32'd299, 32'd92, 32'd5105, 32'd18671},
{32'd13119, -32'd4424, 32'd4611, -32'd8834},
{32'd4328, -32'd9376, 32'd7228, -32'd7727},
{32'd304, 32'd3517, -32'd4039, 32'd6237},
{-32'd7516, -32'd1077, 32'd729, -32'd3730},
{-32'd3415, -32'd2683, 32'd7140, 32'd9199},
{32'd58, -32'd1641, -32'd7322, 32'd2918},
{-32'd6187, 32'd1036, -32'd9154, -32'd6625},
{32'd1485, -32'd4115, -32'd1443, 32'd15879},
{-32'd7273, -32'd4762, -32'd6548, -32'd1240},
{-32'd11297, -32'd5518, -32'd7799, -32'd9122},
{32'd13072, 32'd1441, 32'd1374, -32'd11505},
{-32'd17223, 32'd146, -32'd2559, -32'd3153},
{-32'd1475, -32'd4874, -32'd11244, 32'd4816},
{-32'd478, -32'd6685, -32'd8489, -32'd2160},
{32'd786, -32'd6014, -32'd5863, -32'd7141},
{32'd5317, 32'd5166, -32'd1004, 32'd2786},
{32'd667, -32'd132, 32'd13350, 32'd13594},
{-32'd10169, -32'd18, -32'd2131, -32'd9046},
{-32'd15828, -32'd3248, 32'd7021, 32'd9323},
{-32'd9457, -32'd954, 32'd3268, -32'd4938},
{32'd5248, -32'd602, 32'd7322, -32'd8244},
{32'd12461, -32'd2347, -32'd5502, -32'd3370},
{-32'd2378, -32'd4174, 32'd30, 32'd5371},
{-32'd8726, 32'd2708, -32'd4414, 32'd2205},
{32'd4545, -32'd6138, -32'd46, 32'd4172},
{32'd102, 32'd5354, 32'd5817, -32'd3604},
{-32'd2654, -32'd6178, -32'd981, -32'd540},
{-32'd3487, -32'd2010, -32'd3096, -32'd5395},
{-32'd9919, -32'd5219, -32'd6568, -32'd7091},
{-32'd1648, 32'd882, 32'd7029, 32'd6981},
{-32'd6466, 32'd1222, -32'd5620, -32'd3716},
{32'd856, -32'd4755, -32'd5674, 32'd218},
{32'd13674, 32'd9485, -32'd5030, 32'd3397},
{-32'd625, 32'd2939, 32'd2843, -32'd6291},
{32'd5116, -32'd2274, -32'd8758, -32'd4207},
{-32'd1343, 32'd5712, 32'd5130, -32'd6455},
{-32'd4980, 32'd11301, -32'd5590, 32'd13913},
{-32'd3635, -32'd3493, 32'd8112, 32'd6121},
{-32'd4823, -32'd15859, -32'd3040, -32'd5400},
{-32'd9582, 32'd5265, 32'd3659, 32'd154},
{-32'd9236, 32'd52, -32'd9962, -32'd10137},
{32'd6502, 32'd8289, 32'd9820, 32'd10672},
{-32'd4084, -32'd5526, 32'd996, 32'd1167},
{32'd1209, 32'd3604, -32'd2092, 32'd10235},
{32'd3253, 32'd6865, -32'd2543, -32'd1086},
{32'd10758, -32'd5953, -32'd2332, 32'd7568},
{32'd4838, -32'd1122, -32'd6569, -32'd8035},
{32'd11022, 32'd8960, 32'd3015, 32'd4307},
{-32'd11149, -32'd44, -32'd10094, 32'd1682},
{32'd4696, -32'd804, 32'd3662, -32'd5558},
{32'd4241, 32'd3541, 32'd1527, -32'd4487},
{-32'd1313, 32'd1699, -32'd7526, -32'd3866},
{-32'd9351, -32'd308, -32'd4765, -32'd7989},
{-32'd15295, -32'd4840, 32'd2311, -32'd6914},
{-32'd831, 32'd2568, -32'd6542, 32'd1992},
{-32'd3586, 32'd3099, -32'd10873, -32'd1661},
{32'd1840, -32'd4210, 32'd918, 32'd5248},
{32'd745, -32'd8157, -32'd7981, -32'd6453},
{32'd4627, 32'd5052, 32'd4695, -32'd2386},
{-32'd2776, 32'd4076, -32'd10822, -32'd7925},
{32'd4225, -32'd3700, -32'd9404, -32'd5558},
{-32'd5591, 32'd5055, -32'd2856, -32'd8308},
{32'd5304, 32'd9061, -32'd3830, -32'd10328},
{-32'd625, 32'd4964, 32'd2820, 32'd6025},
{-32'd8966, 32'd11913, -32'd3552, -32'd7983},
{-32'd10147, -32'd5628, -32'd7176, -32'd5182},
{-32'd7352, -32'd886, -32'd6691, -32'd7919},
{32'd5331, -32'd4077, 32'd9934, 32'd977},
{-32'd71, -32'd6570, 32'd9088, 32'd8659},
{32'd2773, 32'd168, -32'd6430, -32'd4155},
{32'd5810, 32'd4566, 32'd4324, 32'd4944},
{32'd1190, -32'd3698, 32'd10873, -32'd1975},
{-32'd6604, 32'd6186, 32'd4034, -32'd300},
{-32'd7866, 32'd2404, -32'd1093, 32'd2807},
{32'd1912, -32'd5341, 32'd191, -32'd12583},
{-32'd1911, -32'd6808, -32'd3860, 32'd2236},
{32'd13577, 32'd192, 32'd1828, -32'd1447},
{32'd8085, -32'd11019, -32'd4963, 32'd1201},
{-32'd2034, 32'd3254, 32'd7766, 32'd2797},
{32'd12625, -32'd4651, -32'd209, -32'd3877},
{32'd4983, 32'd4023, 32'd5651, -32'd6877},
{32'd3006, 32'd1168, 32'd13449, -32'd4248},
{32'd4486, -32'd3480, 32'd6431, 32'd7726},
{32'd3275, -32'd4659, -32'd13400, 32'd3458},
{-32'd9684, 32'd6966, 32'd13392, 32'd3135},
{32'd10843, -32'd4786, -32'd7691, -32'd1733},
{32'd17969, -32'd1886, -32'd11168, 32'd5969},
{32'd510, 32'd5581, -32'd8468, -32'd4363},
{-32'd2440, 32'd6922, -32'd2218, -32'd12441},
{-32'd6821, 32'd9194, 32'd634, -32'd12337},
{-32'd2684, -32'd3702, -32'd1066, -32'd10770},
{32'd8419, -32'd4612, -32'd10864, -32'd6402},
{-32'd5580, -32'd9462, -32'd3095, -32'd1266},
{32'd7611, -32'd8562, -32'd6041, 32'd12843},
{-32'd1772, 32'd86, 32'd6780, -32'd5904},
{-32'd3600, 32'd8872, 32'd3352, -32'd4905},
{32'd596, 32'd499, 32'd485, -32'd1112},
{-32'd11579, -32'd539, 32'd285, 32'd3569},
{32'd6312, -32'd1382, -32'd5773, -32'd7736},
{32'd4557, 32'd5297, 32'd3486, -32'd5829},
{-32'd5526, -32'd9953, -32'd15220, -32'd1537},
{32'd966, -32'd6574, -32'd7605, 32'd2041},
{32'd9726, 32'd11646, -32'd804, -32'd809},
{-32'd9041, -32'd110, -32'd11723, -32'd4179},
{-32'd6013, -32'd3200, -32'd9801, -32'd8285},
{-32'd111, -32'd9946, -32'd3752, -32'd971},
{-32'd2336, 32'd452, 32'd2907, 32'd3904},
{32'd12493, 32'd654, -32'd2836, 32'd4180},
{-32'd4969, 32'd2606, -32'd4382, 32'd11635},
{-32'd506, -32'd6283, -32'd7697, -32'd1311},
{-32'd1758, 32'd975, -32'd3175, -32'd11871},
{-32'd632, -32'd14332, -32'd1319, -32'd3930},
{-32'd2727, 32'd4491, -32'd55, 32'd1354},
{-32'd2064, -32'd2868, -32'd4101, -32'd8318},
{32'd9460, 32'd2829, 32'd9459, 32'd4071},
{-32'd5807, 32'd15515, 32'd5312, -32'd2554},
{-32'd3519, -32'd371, 32'd1141, -32'd4462},
{-32'd5147, -32'd7355, 32'd8649, -32'd532},
{32'd2314, -32'd3865, 32'd9228, 32'd1204},
{32'd6362, -32'd1941, -32'd1544, -32'd1947},
{32'd7374, 32'd330, -32'd851, 32'd1884},
{-32'd18118, 32'd5485, -32'd6197, -32'd5783},
{32'd7149, 32'd2007, 32'd7804, -32'd7375},
{32'd10865, 32'd11142, 32'd1672, 32'd4566},
{-32'd10603, -32'd8087, -32'd2816, 32'd4729},
{-32'd9304, 32'd5315, 32'd12547, -32'd2031},
{-32'd3510, -32'd6468, -32'd6810, 32'd3109},
{-32'd4227, 32'd5577, -32'd2017, 32'd958},
{32'd1225, 32'd8060, 32'd749, -32'd8758},
{-32'd1457, -32'd1776, 32'd3069, 32'd1438},
{-32'd3437, -32'd5870, -32'd1799, -32'd184},
{-32'd5950, -32'd7675, -32'd8766, -32'd13726},
{32'd18722, -32'd3159, -32'd7388, 32'd1184},
{32'd779, -32'd1970, 32'd14211, 32'd7378},
{32'd2723, -32'd4736, -32'd6334, 32'd3383},
{32'd4256, 32'd2363, 32'd2961, 32'd1000},
{32'd1635, 32'd1141, -32'd7267, -32'd1886},
{32'd5902, 32'd3601, 32'd5319, -32'd3530},
{32'd11934, 32'd6309, 32'd1908, 32'd13210},
{32'd6867, 32'd1349, -32'd8537, 32'd5014},
{-32'd5348, 32'd1139, -32'd1143, -32'd7679},
{-32'd1659, -32'd3115, -32'd5255, 32'd4682},
{32'd3797, -32'd8660, -32'd11240, 32'd3708},
{-32'd9248, 32'd1, -32'd5947, 32'd9046},
{-32'd8408, -32'd5106, 32'd8603, 32'd1841},
{32'd5613, -32'd3982, 32'd395, -32'd8332},
{-32'd441, 32'd1835, -32'd3812, -32'd3112},
{-32'd6573, 32'd6035, -32'd9634, -32'd1260},
{-32'd4085, 32'd7179, 32'd7369, -32'd2289},
{-32'd464, -32'd1138, -32'd9392, 32'd2284},
{32'd3942, 32'd1957, 32'd1981, -32'd8622},
{-32'd6885, -32'd8943, -32'd7179, 32'd1874},
{-32'd2554, 32'd600, -32'd5652, -32'd738},
{32'd3149, -32'd2222, 32'd5438, 32'd6213},
{32'd754, 32'd6918, 32'd1364, 32'd6409},
{32'd10142, -32'd9012, 32'd4297, 32'd498},
{-32'd4737, 32'd88, -32'd2371, -32'd4386},
{-32'd1429, 32'd5025, -32'd627, 32'd4371},
{-32'd5627, -32'd3350, -32'd529, 32'd2692},
{-32'd3263, -32'd5692, 32'd1368, -32'd8289},
{-32'd2516, 32'd242, -32'd604, -32'd3701},
{-32'd11591, 32'd7463, -32'd4648, 32'd2737},
{32'd1320, 32'd1043, 32'd5422, -32'd5171},
{-32'd9527, 32'd671, 32'd13752, -32'd10602},
{-32'd2979, 32'd7883, 32'd3113, -32'd5937},
{-32'd802, -32'd1537, -32'd2529, -32'd971},
{-32'd7807, -32'd6749, -32'd7982, 32'd11309},
{32'd388, 32'd3356, 32'd538, -32'd6119},
{32'd2930, -32'd4137, 32'd4182, -32'd10},
{-32'd10318, 32'd3995, -32'd2340, -32'd7525},
{-32'd8912, 32'd103, 32'd2801, -32'd3226},
{32'd622, -32'd7831, -32'd10650, 32'd4697},
{-32'd8100, 32'd4373, 32'd6621, -32'd3663},
{32'd7385, -32'd5550, 32'd3500, 32'd8460},
{32'd223, 32'd7285, 32'd2072, 32'd3286},
{-32'd4553, 32'd468, -32'd6755, 32'd2687},
{-32'd1396, 32'd5828, -32'd222, 32'd9668},
{-32'd4281, -32'd2158, 32'd6728, 32'd348},
{32'd11455, -32'd2230, -32'd737, -32'd8097},
{32'd10781, -32'd5601, 32'd7618, 32'd3991},
{-32'd99, -32'd80, 32'd3408, 32'd7854},
{-32'd19461, 32'd3225, -32'd11897, -32'd772},
{-32'd12911, 32'd305, 32'd1906, -32'd1861},
{-32'd7361, -32'd4647, -32'd158, -32'd7589},
{-32'd5945, -32'd4565, -32'd10733, -32'd521},
{32'd96, -32'd2357, 32'd539, -32'd3211},
{-32'd4960, 32'd2227, -32'd2743, 32'd160},
{-32'd6605, 32'd5064, -32'd1261, -32'd5859},
{-32'd13509, -32'd3664, -32'd2242, 32'd13806},
{32'd11000, 32'd4933, 32'd2645, -32'd6294},
{-32'd6617, -32'd3205, -32'd9242, -32'd5456},
{-32'd2754, -32'd1144, -32'd5959, 32'd773},
{32'd15235, -32'd1093, -32'd4205, -32'd4680},
{-32'd10311, -32'd14451, -32'd12554, -32'd5807},
{32'd1785, 32'd4018, 32'd5129, -32'd6433},
{32'd994, 32'd9650, 32'd3755, 32'd1233},
{-32'd6148, -32'd1436, -32'd14723, 32'd6246},
{32'd994, -32'd5689, -32'd2557, -32'd8957},
{-32'd1667, 32'd243, 32'd3713, -32'd2529},
{32'd1410, -32'd10889, 32'd8737, 32'd5205},
{32'd10291, 32'd732, -32'd3435, -32'd6462},
{-32'd3660, 32'd1835, -32'd7691, 32'd4271},
{-32'd4012, -32'd7391, -32'd13309, 32'd6171},
{32'd1831, 32'd6236, 32'd1603, -32'd586},
{-32'd7730, 32'd1843, 32'd3078, 32'd8625},
{32'd8371, -32'd3293, -32'd7223, 32'd4728},
{-32'd10892, 32'd1098, -32'd3605, 32'd5305},
{-32'd6900, -32'd710, -32'd6172, 32'd115},
{32'd3297, 32'd3777, 32'd5509, -32'd4982},
{32'd2714, 32'd600, -32'd6151, 32'd2553},
{-32'd5082, 32'd1446, 32'd6327, -32'd20384},
{-32'd7705, 32'd805, 32'd978, 32'd5419},
{-32'd7019, 32'd2391, -32'd1240, -32'd1772},
{-32'd3798, -32'd1654, 32'd3024, 32'd2056},
{32'd2033, -32'd3935, -32'd1479, -32'd3078},
{-32'd10745, -32'd2005, 32'd2923, 32'd10509},
{32'd9588, -32'd3199, -32'd3389, -32'd8706},
{32'd9434, -32'd5352, 32'd897, 32'd441},
{-32'd500, -32'd2503, 32'd3414, -32'd5144},
{-32'd9938, -32'd2787, -32'd3060, 32'd11007},
{-32'd2699, -32'd8422, -32'd9596, 32'd7240},
{32'd1782, 32'd6639, 32'd5827, 32'd1211},
{-32'd4999, -32'd3587, 32'd20857, 32'd2016},
{32'd1008, -32'd3596, -32'd2807, 32'd12367},
{-32'd2204, -32'd1147, -32'd7278, -32'd6456},
{-32'd382, -32'd5191, 32'd4301, 32'd395},
{32'd5919, -32'd4565, 32'd2305, -32'd6052},
{32'd3553, 32'd11499, 32'd9025, 32'd778},
{-32'd345, -32'd8251, 32'd7554, -32'd7313},
{-32'd166, -32'd8046, -32'd9835, -32'd4812},
{32'd7376, -32'd7018, -32'd9712, 32'd2745},
{32'd2730, -32'd709, 32'd1511, -32'd10930},
{32'd13928, 32'd5436, 32'd8354, -32'd2087},
{32'd16254, -32'd5388, -32'd3041, -32'd3554},
{32'd17123, -32'd1381, 32'd8014, -32'd1242},
{-32'd1388, 32'd720, 32'd8941, 32'd2583},
{-32'd1030, -32'd3561, -32'd5807, 32'd4388},
{32'd5711, -32'd2315, 32'd2427, -32'd1261},
{32'd812, -32'd5775, -32'd1923, -32'd3835},
{-32'd2345, -32'd1214, -32'd1145, -32'd3241},
{-32'd4793, 32'd6705, -32'd9483, 32'd3208},
{-32'd12620, -32'd4735, 32'd797, 32'd6563},
{-32'd3707, 32'd6391, 32'd3903, -32'd2145},
{32'd3785, -32'd1447, -32'd7404, -32'd8726},
{32'd6958, 32'd7662, 32'd5932, -32'd1730},
{-32'd16730, 32'd524, 32'd1418, 32'd1101},
{-32'd8832, -32'd3902, -32'd7324, 32'd10888},
{32'd10078, -32'd5230, -32'd7237, 32'd553},
{32'd1427, 32'd4503, 32'd3440, -32'd248},
{32'd8697, 32'd4054, 32'd12693, 32'd9533},
{32'd2371, 32'd2858, 32'd274, 32'd6367}
},
{{-32'd7218, 32'd2973, -32'd18139, 32'd3540},
{-32'd12615, 32'd6049, -32'd8331, 32'd3388},
{32'd8534, 32'd6389, 32'd3472, -32'd3223},
{-32'd3513, -32'd3581, 32'd7201, -32'd4284},
{32'd5573, 32'd13891, -32'd117, 32'd3355},
{32'd7917, 32'd2993, -32'd1207, -32'd4741},
{32'd14031, 32'd804, 32'd3042, -32'd10292},
{-32'd7103, -32'd811, 32'd419, -32'd3110},
{32'd15478, 32'd3817, 32'd6336, -32'd239},
{32'd4642, 32'd3757, 32'd9055, -32'd4567},
{32'd15786, -32'd9930, 32'd8628, -32'd5483},
{-32'd5882, 32'd1789, -32'd930, -32'd12260},
{32'd5139, -32'd1075, 32'd8124, 32'd8697},
{-32'd9427, -32'd19480, -32'd4591, 32'd679},
{32'd2350, -32'd18033, 32'd7470, 32'd7324},
{-32'd214, 32'd672, 32'd5201, 32'd9364},
{32'd19960, -32'd7287, -32'd13280, 32'd4469},
{-32'd9481, -32'd4932, 32'd1312, 32'd555},
{-32'd13741, -32'd8150, -32'd1905, -32'd9098},
{32'd7269, 32'd13039, -32'd7959, 32'd1980},
{32'd6825, 32'd10906, -32'd2701, 32'd9185},
{-32'd1322, 32'd90, -32'd8229, 32'd4858},
{32'd4289, -32'd3708, -32'd7854, 32'd9948},
{32'd3420, -32'd11886, -32'd9157, -32'd222},
{32'd10738, 32'd9751, 32'd1457, -32'd7636},
{-32'd10712, -32'd1407, -32'd2560, 32'd3903},
{-32'd4976, -32'd6283, 32'd3484, 32'd3161},
{32'd4328, 32'd1963, 32'd1330, 32'd2274},
{32'd4675, 32'd2050, -32'd5989, -32'd970},
{-32'd9961, 32'd699, 32'd3390, 32'd3512},
{32'd5548, 32'd3233, -32'd13117, 32'd11660},
{32'd1776, -32'd1616, -32'd5970, -32'd5159},
{-32'd3835, 32'd6734, 32'd4045, -32'd7643},
{-32'd12087, 32'd3834, -32'd5863, 32'd4516},
{32'd9172, -32'd2260, 32'd6729, -32'd10791},
{32'd6562, 32'd3458, 32'd11399, -32'd4028},
{-32'd5915, 32'd5836, -32'd6083, -32'd5980},
{32'd654, -32'd4087, -32'd446, 32'd375},
{32'd11892, -32'd1400, -32'd10969, 32'd3936},
{-32'd9053, -32'd18047, 32'd8533, -32'd2709},
{32'd10683, 32'd9112, 32'd4013, -32'd10630},
{32'd12560, -32'd4656, 32'd8716, -32'd709},
{32'd1994, -32'd18989, -32'd6981, -32'd11284},
{-32'd10185, -32'd13079, -32'd474, 32'd4961},
{-32'd11189, -32'd1837, -32'd9794, -32'd387},
{32'd2878, -32'd6329, -32'd2607, -32'd3228},
{32'd11337, 32'd7778, 32'd426, 32'd471},
{-32'd15432, -32'd5217, -32'd9263, 32'd6498},
{32'd2832, -32'd10804, 32'd4718, -32'd2731},
{-32'd8500, -32'd2479, -32'd5704, -32'd638},
{-32'd3318, 32'd7747, -32'd7361, 32'd8495},
{-32'd2262, -32'd5277, 32'd9738, -32'd12540},
{32'd6823, -32'd2808, -32'd18058, -32'd9300},
{-32'd1042, 32'd525, 32'd1647, 32'd3920},
{32'd8485, 32'd7188, 32'd15541, -32'd4759},
{-32'd3628, -32'd7651, -32'd11005, 32'd20069},
{-32'd1173, -32'd4723, -32'd2540, 32'd1174},
{-32'd7941, -32'd3206, 32'd1023, 32'd8760},
{-32'd9505, -32'd11598, -32'd293, -32'd7792},
{-32'd6497, -32'd12431, -32'd8031, -32'd6518},
{-32'd10604, 32'd16104, -32'd6196, 32'd12245},
{32'd7258, -32'd6557, 32'd7272, -32'd15460},
{-32'd569, -32'd354, -32'd3042, 32'd3735},
{-32'd1033, -32'd8226, 32'd2776, 32'd5782},
{-32'd2145, 32'd3833, 32'd1715, -32'd5584},
{-32'd2365, -32'd4714, 32'd5332, -32'd3425},
{-32'd7639, 32'd10001, -32'd17626, 32'd6894},
{32'd1403, 32'd7323, -32'd7050, -32'd3967},
{-32'd7792, 32'd6668, 32'd1657, -32'd2518},
{-32'd722, 32'd3554, 32'd2375, -32'd6382},
{32'd731, 32'd3813, -32'd10752, -32'd1044},
{-32'd4170, -32'd10307, -32'd6152, 32'd3455},
{32'd3390, -32'd12674, -32'd2260, 32'd5896},
{-32'd5924, 32'd163, 32'd991, 32'd7000},
{32'd695, -32'd2055, -32'd1226, -32'd5510},
{32'd125, 32'd21147, 32'd4023, 32'd7124},
{-32'd10540, -32'd8, -32'd4722, 32'd5913},
{32'd4617, -32'd11418, -32'd4365, 32'd2557},
{32'd1159, 32'd227, 32'd3887, 32'd2737},
{-32'd3974, 32'd1193, 32'd6129, 32'd1946},
{-32'd5372, 32'd9825, 32'd2226, -32'd17981},
{-32'd2286, -32'd4048, 32'd3327, -32'd10657},
{-32'd150, 32'd6972, -32'd1627, -32'd669},
{32'd13474, 32'd8390, -32'd15171, -32'd9515},
{-32'd11463, -32'd569, -32'd4601, 32'd1943},
{32'd2875, -32'd11129, -32'd9356, 32'd16485},
{32'd13333, 32'd9258, -32'd2113, -32'd5750},
{-32'd2845, -32'd9644, -32'd563, 32'd5074},
{32'd237, 32'd5566, -32'd1553, 32'd6529},
{-32'd3037, 32'd1703, -32'd17486, -32'd5039},
{32'd6383, 32'd3208, 32'd3525, -32'd14956},
{-32'd3718, -32'd103, -32'd1818, 32'd13629},
{-32'd3689, -32'd955, 32'd6690, -32'd9490},
{32'd7833, 32'd3389, 32'd1145, -32'd5185},
{32'd2244, 32'd7563, -32'd2001, -32'd763},
{32'd2763, 32'd15795, -32'd12061, -32'd696},
{32'd7624, -32'd9126, 32'd3326, -32'd7491},
{-32'd657, 32'd3330, 32'd1623, 32'd2387},
{32'd7332, 32'd10386, 32'd1538, -32'd20107},
{32'd21, -32'd6816, 32'd2323, -32'd4896},
{-32'd9697, 32'd2433, -32'd16472, -32'd6970},
{32'd12195, 32'd5366, -32'd7071, -32'd8213},
{32'd4530, 32'd40, 32'd1213, -32'd4742},
{32'd15587, -32'd5021, -32'd7300, -32'd2839},
{32'd6949, -32'd4783, -32'd2473, -32'd1718},
{32'd5672, -32'd478, 32'd3620, -32'd3837},
{32'd5063, -32'd2461, 32'd2898, 32'd5284},
{32'd8227, -32'd2856, -32'd2531, 32'd16116},
{32'd3291, 32'd3834, -32'd11063, -32'd4060},
{-32'd4804, -32'd2481, -32'd20277, 32'd1083},
{32'd2103, 32'd4465, -32'd3000, -32'd8003},
{32'd3420, 32'd4889, 32'd2935, -32'd13242},
{32'd20277, 32'd1667, 32'd1108, -32'd5926},
{32'd689, 32'd3315, 32'd5721, -32'd19229},
{-32'd4536, -32'd3778, -32'd9069, -32'd351},
{32'd4069, -32'd5759, -32'd6084, -32'd2062},
{32'd7144, -32'd11111, -32'd10743, -32'd12376},
{32'd3504, -32'd860, 32'd10066, 32'd5657},
{32'd3264, -32'd13598, 32'd3093, 32'd5435},
{32'd6710, -32'd9208, 32'd7181, 32'd10065},
{32'd665, 32'd7557, 32'd7347, -32'd159},
{-32'd7907, 32'd353, 32'd11698, 32'd5076},
{-32'd13102, -32'd1298, 32'd6056, 32'd4663},
{32'd6160, 32'd2261, -32'd8924, -32'd16586},
{32'd6619, -32'd4102, -32'd4469, -32'd306},
{32'd12037, 32'd12491, -32'd8924, -32'd351},
{-32'd1968, -32'd9368, 32'd12436, -32'd11173},
{-32'd4865, -32'd5607, 32'd4330, -32'd3011},
{32'd4303, 32'd166, -32'd7418, -32'd1464},
{32'd3631, 32'd14533, -32'd7095, 32'd13389},
{32'd4009, 32'd2108, 32'd2413, -32'd2199},
{32'd2534, 32'd15799, 32'd3948, -32'd11465},
{-32'd382, 32'd4263, -32'd18981, -32'd5374},
{32'd3308, 32'd168, 32'd6570, -32'd3167},
{32'd4794, 32'd11646, 32'd4971, -32'd9810},
{32'd4152, -32'd10987, -32'd1919, 32'd2017},
{-32'd12771, 32'd9194, -32'd2711, 32'd1338},
{32'd9291, 32'd5730, -32'd16474, -32'd3280},
{32'd7835, -32'd310, 32'd1522, 32'd5319},
{-32'd20044, -32'd6458, 32'd7546, -32'd4470},
{32'd9195, 32'd2733, -32'd4386, 32'd5283},
{32'd5380, -32'd11548, -32'd6701, 32'd9203},
{32'd1554, -32'd3847, 32'd1154, 32'd14878},
{32'd7373, -32'd1567, 32'd457, -32'd10822},
{-32'd2615, 32'd8730, -32'd12962, 32'd3341},
{32'd827, -32'd4736, 32'd9625, 32'd11224},
{-32'd6538, -32'd8973, -32'd13284, 32'd4651},
{-32'd6510, -32'd12025, -32'd2979, -32'd8746},
{32'd4755, 32'd15956, 32'd6029, 32'd8693},
{-32'd13175, -32'd14620, -32'd6505, -32'd4728},
{32'd645, -32'd338, -32'd9254, 32'd6200},
{32'd8275, 32'd16502, 32'd10040, -32'd3754},
{-32'd895, -32'd14101, -32'd11442, 32'd5767},
{32'd865, -32'd4434, -32'd9639, 32'd8679},
{32'd7044, -32'd2013, -32'd9927, 32'd440},
{-32'd5722, -32'd1560, 32'd10411, -32'd10045},
{32'd975, 32'd2527, 32'd1214, -32'd5413},
{32'd11493, -32'd2206, -32'd3684, -32'd13476},
{32'd1848, -32'd9459, -32'd6313, 32'd1333},
{-32'd9295, -32'd1902, 32'd8431, -32'd14565},
{32'd5543, 32'd4371, 32'd12319, -32'd7959},
{-32'd20222, 32'd11959, 32'd6200, -32'd4470},
{32'd15741, -32'd4766, -32'd4505, -32'd4241},
{32'd493, 32'd492, 32'd2141, -32'd7100},
{32'd7346, 32'd3354, 32'd10787, 32'd11228},
{-32'd4259, 32'd5383, -32'd29, -32'd3718},
{-32'd838, 32'd16711, 32'd4324, 32'd4059},
{32'd7758, 32'd609, -32'd3492, 32'd2162},
{-32'd4240, -32'd3600, -32'd12786, -32'd4246},
{-32'd5286, -32'd4258, 32'd3316, 32'd6067},
{-32'd4958, -32'd10864, 32'd1808, -32'd3873},
{-32'd6322, 32'd18888, -32'd7967, -32'd5214},
{32'd2482, 32'd325, -32'd1387, -32'd9541},
{-32'd3591, 32'd4364, 32'd13841, -32'd3323},
{-32'd5734, -32'd4059, 32'd7147, 32'd12721},
{-32'd867, 32'd3859, -32'd2705, 32'd9192},
{-32'd4845, 32'd14928, -32'd2437, -32'd3229},
{-32'd5106, 32'd3206, 32'd5765, 32'd10525},
{32'd3966, -32'd140, 32'd4975, 32'd3675},
{-32'd10957, -32'd7165, -32'd12835, 32'd3569},
{-32'd8633, 32'd2706, -32'd1173, 32'd8061},
{-32'd1083, 32'd788, -32'd1219, -32'd7062},
{-32'd5329, 32'd11822, -32'd7825, 32'd4513},
{-32'd2621, -32'd6697, -32'd14041, -32'd1392},
{32'd7746, 32'd8279, -32'd1395, -32'd3733},
{32'd8107, 32'd1288, 32'd4593, -32'd4232},
{32'd14660, 32'd62, 32'd2848, -32'd8530},
{32'd8926, -32'd577, 32'd14742, -32'd455},
{-32'd9477, -32'd1161, 32'd3068, 32'd8881},
{-32'd13439, -32'd7452, 32'd3704, 32'd3303},
{-32'd1313, 32'd8245, 32'd12000, -32'd7563},
{-32'd3299, -32'd10144, 32'd5256, -32'd6305},
{32'd8686, 32'd773, 32'd1692, 32'd5590},
{32'd250, -32'd7099, -32'd139, 32'd830},
{-32'd869, 32'd4972, 32'd2250, 32'd9419},
{32'd6746, -32'd12584, -32'd9624, -32'd931},
{-32'd6302, -32'd4669, -32'd10263, 32'd12079},
{-32'd2517, -32'd5703, -32'd4732, 32'd11993},
{-32'd12058, -32'd1820, -32'd13112, -32'd274},
{32'd4707, 32'd5634, 32'd4242, -32'd12208},
{-32'd9435, 32'd1165, -32'd3555, 32'd1138},
{32'd7322, 32'd1496, -32'd13007, 32'd9899},
{-32'd881, -32'd3858, -32'd4848, -32'd1400},
{32'd7992, 32'd3829, -32'd4944, 32'd4380},
{32'd5940, 32'd5566, -32'd5023, -32'd1525},
{-32'd8227, -32'd6826, -32'd6853, -32'd6001},
{-32'd563, 32'd2428, 32'd3147, -32'd5364},
{-32'd7115, -32'd7069, -32'd10147, 32'd24146},
{-32'd4786, 32'd8459, -32'd369, 32'd5688},
{-32'd1027, 32'd10083, -32'd9861, -32'd17129},
{32'd1277, 32'd3182, -32'd7373, 32'd5916},
{32'd8722, -32'd1936, -32'd5811, 32'd11240},
{-32'd4102, 32'd1902, 32'd3896, 32'd2069},
{-32'd5462, -32'd4799, 32'd4010, 32'd45},
{-32'd11955, -32'd9324, -32'd9325, 32'd3928},
{-32'd5484, -32'd4369, 32'd1025, 32'd7520},
{32'd1783, -32'd1586, -32'd5867, -32'd1509},
{-32'd116, 32'd2695, -32'd1717, 32'd8396},
{-32'd2272, 32'd2148, -32'd8058, 32'd12377},
{32'd2103, -32'd9019, 32'd10352, 32'd4212},
{32'd6390, -32'd7526, -32'd18165, 32'd6288},
{32'd10998, 32'd7223, 32'd6366, -32'd4870},
{32'd8329, 32'd4546, 32'd7688, -32'd5021},
{-32'd1865, -32'd10513, 32'd11077, 32'd5426},
{-32'd9998, -32'd5321, -32'd3124, -32'd10038},
{32'd1424, 32'd421, -32'd5581, -32'd1633},
{-32'd9278, 32'd4102, 32'd2478, 32'd110},
{-32'd9637, -32'd4998, -32'd714, -32'd6585},
{32'd1627, -32'd2685, 32'd1247, -32'd33},
{32'd12703, -32'd4098, -32'd6181, 32'd807},
{-32'd571, -32'd1213, -32'd2894, 32'd4988},
{-32'd8987, -32'd17757, 32'd6301, -32'd9849},
{-32'd4416, -32'd120, 32'd6207, 32'd5722},
{32'd5162, -32'd2437, -32'd1515, -32'd8749},
{-32'd3664, 32'd5011, 32'd9994, 32'd189},
{-32'd1146, 32'd1886, -32'd608, -32'd13643},
{-32'd9316, 32'd8994, 32'd17063, -32'd5218},
{32'd389, -32'd6362, 32'd3983, 32'd10703},
{-32'd7817, 32'd4837, 32'd426, -32'd5423},
{-32'd68, 32'd143, 32'd615, 32'd650},
{32'd2949, -32'd818, 32'd5068, 32'd600},
{-32'd2794, -32'd5959, -32'd10905, 32'd12560},
{-32'd5252, -32'd1007, -32'd792, -32'd1830},
{-32'd6823, -32'd4827, -32'd6504, 32'd7934},
{32'd9781, 32'd7562, 32'd1583, 32'd918},
{-32'd12201, 32'd8745, -32'd8254, 32'd3540},
{-32'd4496, -32'd55, -32'd2492, -32'd10065},
{32'd9507, -32'd7816, -32'd329, -32'd478},
{32'd5891, 32'd8129, -32'd325, -32'd210},
{32'd8699, -32'd2458, -32'd5515, 32'd5784},
{-32'd1961, 32'd620, 32'd703, 32'd11081},
{-32'd5637, -32'd9785, 32'd13501, -32'd13341},
{32'd3792, 32'd15627, 32'd2279, 32'd12393},
{32'd3295, -32'd14699, -32'd2943, 32'd2077},
{32'd3245, -32'd3985, -32'd4672, 32'd8650},
{-32'd2041, -32'd5371, 32'd7246, -32'd1777},
{32'd4657, 32'd13118, -32'd10924, -32'd2396},
{32'd444, 32'd3177, 32'd9126, 32'd4857},
{32'd912, -32'd3023, 32'd1347, -32'd10580},
{32'd1833, -32'd8293, -32'd2485, -32'd12212},
{32'd10864, -32'd6583, 32'd4004, -32'd44},
{32'd2084, 32'd7755, -32'd3151, -32'd1338},
{-32'd5049, 32'd7274, 32'd3767, -32'd3775},
{-32'd9845, -32'd4401, 32'd1419, 32'd9952},
{32'd3682, 32'd11991, -32'd5424, 32'd12080},
{-32'd11915, -32'd117, -32'd1955, 32'd6734},
{-32'd6805, -32'd4860, 32'd13981, -32'd13691},
{32'd1134, 32'd2047, -32'd4940, 32'd4856},
{32'd6103, -32'd12040, 32'd372, -32'd3213},
{-32'd6643, -32'd6828, -32'd11358, 32'd4073},
{32'd4720, 32'd1589, -32'd11616, -32'd807},
{32'd12784, 32'd14169, -32'd7135, -32'd14621},
{32'd5144, -32'd5012, -32'd18831, 32'd8284},
{-32'd6166, -32'd5621, -32'd883, 32'd7131},
{32'd5464, 32'd3733, 32'd1699, -32'd3008},
{-32'd1666, 32'd438, -32'd3309, 32'd3890},
{32'd3651, 32'd1020, 32'd7403, -32'd1088},
{32'd2393, 32'd3914, 32'd3867, 32'd5019},
{-32'd8504, -32'd4187, -32'd2059, -32'd699},
{32'd2284, -32'd8625, -32'd2057, 32'd1994},
{32'd3132, 32'd1682, -32'd3812, -32'd5053},
{32'd9258, 32'd7236, 32'd14748, -32'd10157},
{32'd5602, 32'd2547, 32'd12463, -32'd3889},
{-32'd8129, -32'd5286, -32'd15519, 32'd319},
{32'd11163, 32'd15164, -32'd7336, 32'd19},
{-32'd179, -32'd304, -32'd3851, -32'd6497},
{-32'd7855, -32'd2228, -32'd7380, 32'd1533},
{32'd3104, -32'd8570, -32'd10065, 32'd5113},
{32'd2222, -32'd6539, -32'd1418, 32'd8776},
{32'd5642, -32'd5621, -32'd1584, -32'd23514},
{-32'd4277, -32'd7177, 32'd4819, 32'd212},
{32'd4439, 32'd2685, 32'd8804, -32'd19106},
{-32'd9507, -32'd5373, 32'd8905, -32'd9517},
{-32'd6735, -32'd191, -32'd2110, -32'd6224},
{32'd1152, -32'd5963, 32'd4168, -32'd2309},
{-32'd10573, -32'd374, 32'd312, -32'd1807},
{-32'd4342, 32'd4146, -32'd228, 32'd1627},
{32'd14204, -32'd3634, 32'd3825, -32'd8521},
{32'd4219, 32'd1207, 32'd4353, -32'd1801},
{32'd3103, 32'd3210, 32'd2418, -32'd1415}
},
{{-32'd3838, 32'd8785, 32'd3619, 32'd4724},
{32'd2560, -32'd4905, -32'd6859, 32'd5310},
{-32'd3214, -32'd251, -32'd7445, -32'd5660},
{32'd6056, 32'd6317, -32'd10469, -32'd3687},
{32'd14652, 32'd5632, 32'd2632, -32'd3140},
{-32'd11, -32'd3898, 32'd4781, 32'd4776},
{32'd4962, 32'd8291, 32'd14812, -32'd394},
{-32'd7202, -32'd1568, -32'd10822, 32'd2428},
{-32'd2316, 32'd1881, 32'd1361, 32'd5693},
{32'd5318, 32'd4205, 32'd6259, -32'd440},
{-32'd1199, 32'd1132, 32'd6920, 32'd3948},
{-32'd192, -32'd41, 32'd949, -32'd2822},
{32'd4566, -32'd8386, -32'd144, -32'd13048},
{32'd2064, -32'd339, -32'd5016, 32'd1764},
{32'd1021, -32'd14121, 32'd344, 32'd11762},
{-32'd3174, 32'd3548, 32'd2770, -32'd3499},
{-32'd5186, 32'd13009, 32'd10487, -32'd4897},
{-32'd5878, 32'd12596, -32'd14182, -32'd3372},
{32'd2099, 32'd7352, -32'd9270, 32'd5153},
{32'd9226, -32'd447, 32'd2706, -32'd6614},
{32'd12450, 32'd1731, -32'd2363, 32'd4004},
{-32'd6546, -32'd7463, -32'd7380, -32'd2077},
{32'd5909, 32'd385, 32'd2860, 32'd5413},
{-32'd3409, -32'd2522, -32'd3784, 32'd9096},
{32'd1220, 32'd7567, 32'd5317, -32'd829},
{32'd890, -32'd2546, 32'd4726, 32'd8011},
{-32'd14738, 32'd14005, 32'd5780, 32'd2235},
{32'd4448, 32'd8985, -32'd151, -32'd11516},
{32'd11413, 32'd7505, -32'd2391, -32'd2247},
{32'd99, 32'd5754, -32'd3203, 32'd7851},
{-32'd984, 32'd5524, 32'd13665, 32'd10775},
{-32'd1168, -32'd6072, 32'd2165, 32'd9337},
{-32'd835, 32'd3984, 32'd4896, -32'd2615},
{-32'd5404, -32'd4687, -32'd1849, 32'd929},
{32'd8289, 32'd8235, 32'd8470, -32'd299},
{-32'd2811, 32'd9142, -32'd6973, -32'd107},
{32'd2829, -32'd8057, 32'd7671, 32'd370},
{-32'd2327, -32'd9627, -32'd6086, 32'd11103},
{-32'd4359, -32'd4368, 32'd1834, -32'd4682},
{-32'd12914, 32'd7968, 32'd7625, -32'd5892},
{32'd793, 32'd753, -32'd7695, -32'd12946},
{32'd5531, 32'd11382, -32'd266, -32'd4993},
{-32'd3335, 32'd1247, 32'd10911, -32'd5696},
{-32'd9847, -32'd6030, -32'd10203, -32'd484},
{-32'd16542, -32'd15058, -32'd9535, -32'd9347},
{32'd2378, 32'd2393, 32'd2686, -32'd609},
{32'd3495, -32'd1502, 32'd7151, -32'd2974},
{-32'd16752, -32'd6937, -32'd12447, 32'd3929},
{-32'd4165, 32'd629, 32'd7191, 32'd1836},
{-32'd6877, -32'd4282, 32'd1370, 32'd7120},
{-32'd2250, -32'd10521, -32'd11256, -32'd7819},
{32'd7184, -32'd3104, 32'd6401, 32'd5797},
{32'd5687, 32'd425, -32'd9139, 32'd2329},
{-32'd4783, -32'd11714, -32'd5390, -32'd6066},
{-32'd6997, 32'd16199, -32'd1175, 32'd1720},
{32'd564, -32'd632, 32'd7591, 32'd3202},
{32'd1832, 32'd2523, 32'd4598, -32'd3292},
{-32'd3951, 32'd1389, -32'd5128, 32'd2055},
{-32'd3125, 32'd13277, -32'd9653, 32'd1645},
{32'd6392, -32'd8406, 32'd7037, 32'd7483},
{-32'd4933, 32'd7067, 32'd980, 32'd3511},
{32'd8790, 32'd4912, -32'd4873, -32'd10442},
{-32'd3796, 32'd411, -32'd5480, -32'd5178},
{32'd1805, -32'd6220, -32'd7188, -32'd6669},
{32'd6213, -32'd13867, -32'd9767, 32'd4909},
{32'd11166, 32'd5165, -32'd4683, 32'd2546},
{32'd8773, 32'd1913, 32'd8543, 32'd13110},
{32'd6418, -32'd8711, -32'd1544, 32'd6478},
{-32'd3048, 32'd9579, -32'd10058, -32'd2707},
{32'd12856, -32'd6357, -32'd4364, -32'd2765},
{-32'd5620, 32'd565, 32'd4330, -32'd6875},
{-32'd11067, 32'd6137, 32'd1813, 32'd4038},
{-32'd6848, 32'd6189, -32'd2397, -32'd8505},
{-32'd1028, 32'd6506, 32'd1323, 32'd433},
{32'd5482, 32'd1171, 32'd6931, 32'd9699},
{-32'd3052, 32'd17173, 32'd2249, -32'd7592},
{-32'd12054, -32'd7878, -32'd10035, 32'd3318},
{-32'd1154, 32'd9381, -32'd2372, 32'd11049},
{32'd3436, 32'd2460, 32'd2064, -32'd1036},
{32'd1904, 32'd5496, 32'd3016, 32'd190},
{32'd2543, -32'd1800, -32'd2399, -32'd7648},
{-32'd5882, 32'd1076, -32'd5585, -32'd15994},
{32'd3496, -32'd7225, 32'd4634, 32'd4256},
{32'd7973, -32'd2120, 32'd5894, 32'd6168},
{-32'd13748, 32'd2709, -32'd13652, 32'd379},
{32'd1362, -32'd17605, 32'd2684, -32'd1758},
{32'd7292, 32'd2651, -32'd14609, -32'd6593},
{-32'd10224, -32'd6246, -32'd6597, -32'd2607},
{32'd408, -32'd6064, -32'd5015, 32'd1576},
{32'd3084, 32'd4024, -32'd5025, 32'd8326},
{-32'd110, 32'd3365, 32'd8944, -32'd6434},
{32'd8301, 32'd6733, -32'd9511, 32'd13892},
{-32'd717, 32'd3039, -32'd5766, 32'd527},
{32'd3013, 32'd5731, 32'd8457, 32'd1996},
{-32'd10363, 32'd8316, 32'd1573, 32'd44},
{-32'd2505, 32'd13844, -32'd8936, 32'd3500},
{32'd2827, 32'd2565, 32'd5019, -32'd4876},
{32'd1525, -32'd6002, -32'd6694, -32'd8418},
{-32'd9907, 32'd565, -32'd4895, -32'd9611},
{32'd1788, 32'd9160, -32'd3135, -32'd1442},
{-32'd2776, -32'd14727, 32'd4839, 32'd14453},
{-32'd8884, -32'd3089, 32'd1447, -32'd10307},
{-32'd4270, -32'd12104, 32'd9818, 32'd5834},
{32'd9267, 32'd8001, -32'd340, 32'd8081},
{32'd2294, -32'd2553, 32'd3306, -32'd5503},
{32'd10592, 32'd9298, 32'd15228, 32'd1206},
{32'd1796, -32'd10124, 32'd11524, -32'd5127},
{32'd246, -32'd4951, 32'd4085, -32'd5684},
{32'd1123, 32'd9488, 32'd4026, 32'd5892},
{-32'd10545, -32'd8432, -32'd1430, -32'd853},
{32'd5483, -32'd1266, -32'd5724, -32'd6021},
{-32'd3448, -32'd4595, 32'd384, -32'd7521},
{32'd2842, 32'd6779, 32'd6288, -32'd9706},
{-32'd3687, 32'd12190, -32'd9436, -32'd3812},
{32'd11056, 32'd8947, -32'd4690, 32'd7053},
{32'd5944, 32'd1668, 32'd1407, -32'd1700},
{32'd5161, 32'd4141, 32'd7139, 32'd3627},
{32'd11514, 32'd578, 32'd1940, 32'd4305},
{-32'd2586, -32'd4709, 32'd5323, -32'd3010},
{32'd7620, 32'd10640, 32'd11241, 32'd11218},
{32'd5284, 32'd18694, -32'd14402, 32'd3476},
{32'd6904, 32'd1859, -32'd10503, 32'd255},
{-32'd1206, -32'd245, -32'd6059, 32'd2722},
{32'd13561, 32'd1949, 32'd4510, -32'd3906},
{-32'd4654, -32'd3732, -32'd16601, 32'd2158},
{-32'd3776, 32'd3897, 32'd5739, 32'd110},
{-32'd4642, -32'd54, -32'd6125, -32'd6172},
{32'd386, -32'd894, -32'd4399, 32'd1816},
{-32'd1472, -32'd5622, -32'd640, 32'd8528},
{-32'd10557, -32'd7240, 32'd1469, -32'd4043},
{-32'd1000, -32'd485, -32'd2964, -32'd18142},
{-32'd5767, -32'd9619, 32'd5368, -32'd1801},
{-32'd4203, -32'd17154, -32'd305, 32'd3135},
{-32'd12453, -32'd2482, 32'd6675, -32'd4995},
{-32'd1170, -32'd1157, -32'd7148, -32'd4204},
{-32'd15119, -32'd5067, -32'd3467, -32'd10291},
{32'd13582, 32'd742, -32'd9577, -32'd1668},
{-32'd6401, 32'd4732, -32'd1690, -32'd6652},
{32'd11583, 32'd1662, -32'd271, 32'd8426},
{-32'd8582, -32'd10248, -32'd6918, -32'd2939},
{-32'd1166, -32'd6194, 32'd3432, -32'd3470},
{32'd8754, 32'd1245, -32'd6641, -32'd16836},
{32'd4164, 32'd5643, 32'd5254, 32'd9059},
{-32'd5091, -32'd257, 32'd5012, 32'd5304},
{32'd3607, 32'd3216, -32'd2927, 32'd6025},
{-32'd4493, -32'd2465, 32'd6310, -32'd683},
{-32'd12863, -32'd4584, 32'd4996, 32'd13773},
{-32'd16818, 32'd3827, 32'd12458, -32'd857},
{-32'd875, 32'd5020, -32'd3492, -32'd1810},
{-32'd13867, -32'd11424, -32'd5552, 32'd3040},
{-32'd13315, -32'd1636, -32'd8255, 32'd591},
{-32'd3840, 32'd4319, 32'd1066, -32'd5979},
{-32'd2716, -32'd12821, -32'd9605, -32'd6927},
{32'd134, 32'd1460, 32'd9238, -32'd589},
{-32'd6193, -32'd9437, -32'd3455, -32'd2147},
{32'd9969, -32'd14984, -32'd3075, -32'd10199},
{-32'd292, 32'd3009, -32'd3250, -32'd2828},
{32'd4659, 32'd1599, -32'd10072, -32'd5151},
{32'd3356, -32'd10039, -32'd3367, 32'd7195},
{32'd1519, 32'd8829, -32'd1387, -32'd11273},
{-32'd1691, 32'd3385, -32'd6444, -32'd9021},
{32'd2125, 32'd2992, -32'd10912, -32'd5124},
{32'd7203, 32'd2289, 32'd9415, -32'd22760},
{-32'd1439, 32'd2653, 32'd3516, 32'd1336},
{32'd13454, 32'd5271, 32'd21140, -32'd6951},
{32'd2950, -32'd3944, 32'd11068, 32'd5345},
{32'd3544, 32'd3925, 32'd8215, 32'd9621},
{-32'd4829, -32'd4099, -32'd15163, -32'd5884},
{-32'd15596, 32'd4374, 32'd789, -32'd10316},
{-32'd7537, -32'd8776, 32'd2905, 32'd6495},
{-32'd7050, -32'd646, 32'd6, 32'd13929},
{-32'd1340, -32'd1752, -32'd343, 32'd14084},
{32'd7625, 32'd7480, 32'd14340, -32'd3532},
{-32'd7747, -32'd6436, -32'd14048, 32'd4705},
{32'd6292, -32'd6010, 32'd8736, -32'd3590},
{-32'd1962, -32'd2488, -32'd4039, 32'd4322},
{32'd3221, -32'd8449, 32'd150, -32'd1163},
{-32'd2172, 32'd4344, 32'd9059, 32'd5327},
{-32'd1989, 32'd4115, 32'd8082, -32'd6386},
{-32'd20067, -32'd6952, -32'd6948, 32'd13277},
{-32'd12987, -32'd9188, -32'd1299, -32'd3424},
{-32'd6686, -32'd13537, -32'd5879, -32'd1864},
{32'd4717, -32'd151, -32'd853, 32'd3059},
{-32'd5422, -32'd4147, -32'd17149, -32'd7141},
{-32'd174, -32'd2909, -32'd1794, 32'd15024},
{32'd14539, 32'd312, 32'd2603, 32'd3917},
{32'd4752, 32'd3561, -32'd1041, -32'd6558},
{-32'd19117, 32'd7009, -32'd10182, 32'd2175},
{-32'd3938, -32'd9048, 32'd7988, 32'd4937},
{32'd5926, -32'd8466, -32'd5091, -32'd12107},
{32'd362, 32'd8518, -32'd3254, 32'd1874},
{-32'd8991, -32'd3596, 32'd136, -32'd319},
{-32'd3917, -32'd4712, 32'd5761, 32'd20863},
{32'd1480, -32'd5366, -32'd13628, -32'd4915},
{-32'd12509, -32'd7686, -32'd4965, 32'd3227},
{32'd2464, 32'd11973, -32'd134, -32'd9288},
{32'd4196, -32'd1652, 32'd7664, 32'd15163},
{-32'd1955, -32'd1245, 32'd13099, -32'd2414},
{32'd2547, -32'd14570, -32'd9750, -32'd11293},
{32'd4890, 32'd11519, 32'd10640, -32'd17945},
{-32'd4243, -32'd7355, -32'd6089, -32'd3372},
{-32'd3080, 32'd2943, 32'd8149, -32'd2975},
{-32'd7859, 32'd2638, 32'd4332, -32'd7607},
{32'd3866, 32'd6420, 32'd2925, -32'd1535},
{-32'd2756, -32'd1144, -32'd21094, 32'd13683},
{32'd2762, 32'd7155, 32'd358, -32'd3179},
{32'd6811, 32'd6394, 32'd5156, -32'd3202},
{32'd1175, -32'd11689, -32'd2020, 32'd9966},
{-32'd14137, 32'd18424, -32'd193, -32'd8754},
{-32'd8831, 32'd4284, -32'd9739, -32'd3897},
{-32'd6773, 32'd2201, 32'd4079, 32'd6740},
{32'd2792, -32'd5108, 32'd948, 32'd4912},
{32'd2225, -32'd14616, -32'd10696, 32'd3622},
{32'd791, 32'd4747, 32'd5644, 32'd11122},
{-32'd5436, -32'd2531, 32'd3034, 32'd2806},
{-32'd1767, 32'd8647, -32'd9298, 32'd4273},
{32'd36, 32'd6074, -32'd1021, -32'd460},
{-32'd5869, -32'd7736, -32'd5652, 32'd19304},
{-32'd4769, -32'd3863, 32'd12280, 32'd398},
{-32'd2115, 32'd1285, -32'd2382, -32'd6665},
{32'd2969, 32'd3398, 32'd11069, 32'd2640},
{32'd2945, -32'd2951, -32'd2816, 32'd1359},
{-32'd669, -32'd1072, 32'd4110, -32'd3606},
{-32'd4051, 32'd12048, 32'd9575, -32'd5672},
{32'd8229, -32'd10951, -32'd6241, 32'd6663},
{-32'd8712, -32'd7852, 32'd2225, -32'd8349},
{32'd7001, -32'd14633, -32'd12251, 32'd7839},
{32'd3747, -32'd4751, -32'd17795, 32'd5626},
{32'd8105, -32'd4298, 32'd2074, -32'd15502},
{32'd4999, 32'd5106, -32'd1099, -32'd10873},
{-32'd317, 32'd4152, 32'd2643, -32'd899},
{32'd1177, 32'd10632, 32'd1557, -32'd7885},
{32'd3489, 32'd8160, 32'd4676, 32'd10385},
{32'd1008, 32'd2213, -32'd11953, -32'd5956},
{-32'd3434, 32'd6362, -32'd8573, -32'd2313},
{-32'd7815, -32'd741, -32'd17302, 32'd5582},
{32'd8685, -32'd17825, -32'd10315, 32'd675},
{-32'd4959, -32'd3022, 32'd16872, 32'd5093},
{32'd10520, 32'd8115, 32'd10892, 32'd580},
{-32'd247, 32'd21544, -32'd8009, 32'd2957},
{-32'd1856, 32'd9918, 32'd4744, -32'd4128},
{-32'd6077, 32'd11523, -32'd10788, 32'd103},
{-32'd8090, 32'd1009, -32'd2601, 32'd4533},
{32'd3764, -32'd3885, 32'd13520, 32'd19608},
{32'd7438, 32'd4404, 32'd1559, -32'd300},
{32'd2417, 32'd6497, 32'd1757, 32'd7341},
{-32'd5936, -32'd9502, -32'd5694, -32'd3},
{32'd11312, -32'd2829, 32'd7056, 32'd3919},
{-32'd819, 32'd8991, 32'd2362, 32'd2014},
{-32'd236, -32'd6499, 32'd7616, 32'd1841},
{32'd1707, -32'd10043, -32'd4285, 32'd3099},
{-32'd1393, 32'd16268, -32'd5866, -32'd8650},
{-32'd7271, 32'd3106, 32'd13484, -32'd5792},
{-32'd716, -32'd7120, 32'd11015, 32'd14343},
{-32'd10718, -32'd8519, 32'd9742, -32'd457},
{32'd251, -32'd1547, 32'd14048, -32'd6141},
{32'd6447, -32'd10919, 32'd12955, 32'd8303},
{32'd198, -32'd5551, 32'd1038, 32'd1269},
{-32'd9003, 32'd1116, -32'd9179, 32'd739},
{-32'd3117, -32'd914, 32'd4661, 32'd1926},
{32'd4634, 32'd4460, 32'd12851, -32'd6642},
{32'd7422, 32'd4369, -32'd7877, 32'd8167},
{32'd12269, -32'd11110, -32'd10529, 32'd12175},
{32'd10388, 32'd14297, -32'd11305, 32'd33},
{32'd8431, 32'd12619, 32'd1975, 32'd15216},
{-32'd10600, 32'd6414, 32'd3008, -32'd13230},
{32'd16601, 32'd6949, -32'd7044, -32'd8317},
{32'd2135, 32'd23807, -32'd20635, -32'd10775},
{-32'd5929, 32'd3092, -32'd2233, 32'd6093},
{32'd4259, -32'd1935, -32'd18302, 32'd4569},
{32'd1441, 32'd11738, 32'd157, 32'd11977},
{32'd8731, -32'd3711, -32'd1271, 32'd10386},
{32'd2103, -32'd8043, 32'd3203, -32'd14070},
{32'd2720, 32'd2579, -32'd6319, 32'd4261},
{-32'd2760, 32'd4774, -32'd5022, 32'd7754},
{-32'd4862, 32'd3767, 32'd2803, 32'd12287},
{32'd9790, 32'd6615, 32'd4015, -32'd281},
{32'd1707, 32'd13122, 32'd5743, 32'd4665},
{-32'd3250, 32'd2215, -32'd5335, 32'd8237},
{32'd7185, -32'd461, 32'd81, 32'd5849},
{32'd10163, -32'd5920, 32'd4445, 32'd8973},
{32'd3331, 32'd1230, -32'd6103, -32'd6250},
{32'd4878, -32'd867, 32'd13993, 32'd2042},
{32'd1121, -32'd9776, 32'd5881, 32'd13673},
{32'd9229, 32'd18276, 32'd13935, -32'd4100},
{-32'd5384, -32'd12449, -32'd8545, -32'd4250},
{32'd16552, 32'd2161, -32'd2999, -32'd3724},
{32'd5361, -32'd7200, -32'd1897, 32'd14996},
{-32'd102, -32'd5180, -32'd7030, 32'd5530},
{-32'd1345, -32'd11635, -32'd2582, -32'd12555},
{-32'd3773, -32'd1869, 32'd10545, -32'd7437},
{32'd5977, 32'd5914, 32'd7256, -32'd1782},
{32'd4421, -32'd9900, 32'd6399, -32'd30},
{32'd10630, 32'd6762, -32'd19686, -32'd7527},
{-32'd3468, -32'd1321, 32'd10215, -32'd1324},
{-32'd10806, 32'd6972, -32'd3919, 32'd10255},
{32'd3052, 32'd378, -32'd303, -32'd2714},
{32'd9801, 32'd3490, -32'd3838, -32'd17931},
{32'd10138, -32'd1863, 32'd17555, -32'd3263},
{-32'd8993, 32'd4083, -32'd8636, -32'd34}
},
{{32'd14754, 32'd5506, 32'd3626, 32'd4795},
{-32'd4499, 32'd2040, 32'd430, 32'd1880},
{32'd988, -32'd1942, 32'd4186, 32'd190},
{-32'd5850, -32'd4486, 32'd8053, 32'd6159},
{-32'd7775, -32'd1772, 32'd10249, 32'd4113},
{-32'd2369, 32'd175, 32'd1261, 32'd4047},
{32'd4602, 32'd10211, -32'd54, -32'd1111},
{-32'd1360, 32'd9337, -32'd4657, -32'd2382},
{32'd3803, 32'd4480, -32'd1450, 32'd317},
{32'd3663, 32'd468, 32'd7618, 32'd4254},
{-32'd6475, -32'd1613, -32'd1564, 32'd7025},
{-32'd1291, 32'd1833, -32'd7113, -32'd1084},
{-32'd3359, 32'd8617, 32'd14816, 32'd3178},
{-32'd2189, -32'd4996, -32'd749, -32'd8521},
{-32'd7946, 32'd6051, -32'd2327, -32'd1612},
{32'd3567, 32'd4791, -32'd5913, -32'd850},
{32'd3911, 32'd9143, 32'd9448, 32'd700},
{32'd10915, -32'd375, 32'd468, -32'd1682},
{32'd2189, 32'd7645, 32'd4764, -32'd2748},
{32'd10463, -32'd5079, 32'd8309, -32'd434},
{32'd4236, -32'd3169, 32'd2204, 32'd135},
{-32'd4777, -32'd3028, -32'd4831, -32'd1038},
{-32'd710, 32'd814, -32'd956, -32'd3964},
{-32'd5128, -32'd936, -32'd3786, -32'd3548},
{32'd8406, -32'd9018, 32'd1375, 32'd6056},
{-32'd11157, 32'd5957, 32'd5726, 32'd3642},
{-32'd3912, 32'd9233, -32'd1754, -32'd6958},
{32'd8949, 32'd286, 32'd4990, 32'd5806},
{32'd12927, -32'd12257, 32'd3804, 32'd3209},
{-32'd6588, -32'd4547, -32'd4600, -32'd5131},
{32'd1490, 32'd450, 32'd12572, 32'd2791},
{32'd5700, -32'd11360, -32'd1088, -32'd4765},
{32'd20698, 32'd18236, 32'd2630, 32'd2075},
{-32'd9417, 32'd4436, 32'd6426, -32'd6228},
{-32'd3851, 32'd3692, 32'd10035, 32'd1579},
{-32'd3593, -32'd3193, 32'd793, 32'd5352},
{-32'd6867, 32'd3187, -32'd5825, 32'd4040},
{-32'd2432, 32'd17888, -32'd3825, -32'd12306},
{32'd9997, 32'd8048, 32'd5249, -32'd6397},
{32'd19400, 32'd5363, 32'd1204, -32'd9026},
{32'd2170, -32'd9001, 32'd2206, 32'd685},
{-32'd1997, 32'd15973, 32'd4113, 32'd4020},
{-32'd3101, 32'd13619, 32'd1156, -32'd744},
{-32'd5349, -32'd4772, -32'd9537, 32'd1499},
{32'd3304, -32'd2579, -32'd6157, -32'd9522},
{-32'd5723, -32'd5924, 32'd1611, -32'd1248},
{32'd8280, 32'd4851, 32'd2258, -32'd3108},
{-32'd4195, -32'd13737, 32'd1022, -32'd6947},
{32'd182, 32'd4827, -32'd2790, -32'd1777},
{-32'd1697, -32'd3643, -32'd10803, -32'd1552},
{32'd6329, -32'd4694, 32'd677, 32'd3669},
{-32'd4298, -32'd33, -32'd4749, -32'd2889},
{32'd5086, -32'd3504, -32'd3240, -32'd1703},
{-32'd5956, 32'd252, -32'd7515, -32'd3309},
{32'd1330, -32'd2973, -32'd8844, -32'd2045},
{-32'd4117, -32'd11208, 32'd481, -32'd817},
{32'd16337, 32'd17031, 32'd22, -32'd1570},
{32'd1900, 32'd3146, -32'd941, 32'd2353},
{-32'd4895, -32'd8008, -32'd12095, -32'd5720},
{32'd6437, -32'd4370, 32'd6397, 32'd2224},
{32'd2575, 32'd6862, 32'd1803, 32'd2649},
{-32'd13296, -32'd5912, 32'd202, -32'd999},
{-32'd6746, -32'd4445, 32'd1011, -32'd6488},
{-32'd6235, -32'd5817, -32'd4830, 32'd6351},
{-32'd592, 32'd2948, -32'd8655, 32'd1040},
{32'd5234, 32'd2913, 32'd10211, 32'd6516},
{32'd4210, 32'd5266, 32'd1143, -32'd4996},
{-32'd3447, 32'd2589, -32'd1403, -32'd2935},
{32'd7466, -32'd12927, 32'd2493, -32'd2044},
{32'd809, 32'd5351, 32'd3884, 32'd8616},
{32'd3534, -32'd11093, -32'd3300, 32'd1218},
{-32'd6120, 32'd1567, 32'd324, 32'd4465},
{32'd5243, -32'd1200, -32'd2869, 32'd908},
{32'd12795, 32'd12332, 32'd5802, 32'd5489},
{32'd15976, -32'd2174, 32'd2544, 32'd5126},
{-32'd5141, 32'd4664, -32'd3712, -32'd593},
{32'd1156, -32'd12859, -32'd9776, -32'd3948},
{32'd2760, -32'd2219, -32'd4348, 32'd2483},
{-32'd6427, 32'd697, 32'd11072, -32'd1515},
{-32'd5801, -32'd1194, -32'd2992, 32'd3781},
{32'd4581, -32'd11414, -32'd2581, -32'd2071},
{32'd12553, 32'd8110, 32'd683, -32'd2469},
{32'd472, -32'd10874, -32'd846, -32'd457},
{-32'd1141, 32'd6493, -32'd10804, -32'd2063},
{32'd1251, -32'd10286, -32'd1040, -32'd7889},
{32'd5684, 32'd8291, 32'd2521, -32'd987},
{-32'd4722, -32'd77, 32'd5158, -32'd161},
{-32'd9874, 32'd5487, -32'd3478, 32'd208},
{-32'd9084, -32'd655, -32'd319, 32'd3358},
{-32'd12589, -32'd3453, -32'd10327, -32'd7881},
{32'd7607, 32'd12216, 32'd5266, 32'd97},
{32'd1446, 32'd3294, -32'd3276, -32'd125},
{-32'd1757, -32'd1075, 32'd11626, -32'd1438},
{32'd3458, 32'd7014, 32'd7254, -32'd455},
{-32'd9595, -32'd4200, 32'd5543, 32'd1413},
{-32'd31, -32'd2413, -32'd9012, 32'd1161},
{-32'd1906, 32'd10089, 32'd8620, 32'd8},
{-32'd828, 32'd12542, 32'd778, -32'd1466},
{32'd3908, -32'd172, 32'd487, 32'd918},
{-32'd1657, -32'd185, 32'd6843, -32'd790},
{-32'd19479, -32'd7959, -32'd8706, -32'd159},
{-32'd1024, -32'd3008, 32'd2068, -32'd2769},
{-32'd7205, -32'd5455, -32'd445, -32'd4197},
{-32'd7946, -32'd1948, -32'd6074, 32'd10248},
{32'd7140, 32'd470, 32'd10010, 32'd13116},
{32'd524, -32'd12676, -32'd10802, -32'd3356},
{-32'd46, -32'd582, -32'd3623, -32'd5228},
{-32'd13712, -32'd2573, 32'd4461, -32'd7426},
{32'd4289, -32'd1812, 32'd5914, 32'd2544},
{32'd7032, 32'd5044, -32'd11820, 32'd2718},
{-32'd12844, -32'd7912, -32'd2635, 32'd2239},
{32'd11584, -32'd10125, -32'd9144, -32'd855},
{32'd2188, -32'd2044, 32'd2172, 32'd3465},
{-32'd6158, 32'd5974, 32'd5036, 32'd6063},
{-32'd11376, -32'd10449, -32'd10910, -32'd1924},
{32'd4579, -32'd6529, -32'd1389, 32'd5825},
{-32'd14526, -32'd16182, -32'd724, -32'd923},
{32'd73, 32'd1383, -32'd10314, -32'd632},
{32'd5261, -32'd9949, -32'd11813, 32'd811},
{32'd4192, 32'd2436, 32'd10271, 32'd6929},
{-32'd5911, -32'd4196, 32'd3225, -32'd2211},
{-32'd5877, 32'd1887, -32'd1250, 32'd5429},
{32'd12569, -32'd2813, 32'd1880, -32'd1600},
{-32'd3278, -32'd11133, 32'd8360, 32'd1628},
{32'd1762, -32'd8370, 32'd4465, -32'd627},
{32'd3913, 32'd2691, 32'd712, -32'd1364},
{-32'd2600, -32'd8827, -32'd95, -32'd2481},
{-32'd3071, -32'd9923, -32'd808, 32'd8201},
{-32'd4785, 32'd4117, -32'd1625, 32'd654},
{32'd10486, 32'd216, 32'd4782, 32'd9671},
{-32'd1183, 32'd6099, 32'd3436, 32'd2936},
{32'd1383, 32'd335, -32'd386, -32'd4095},
{32'd6848, -32'd14483, -32'd520, 32'd4776},
{32'd4543, -32'd4900, 32'd1539, 32'd912},
{32'd8460, -32'd4545, 32'd136, 32'd8849},
{32'd8605, 32'd1540, -32'd4180, -32'd860},
{-32'd3758, 32'd2682, -32'd21, 32'd2473},
{-32'd8877, -32'd15559, -32'd2003, 32'd2021},
{32'd15253, 32'd2595, 32'd2453, 32'd1376},
{32'd6160, -32'd4131, -32'd1934, -32'd6215},
{32'd9448, 32'd2022, -32'd7076, 32'd5198},
{-32'd2490, -32'd2816, 32'd10432, -32'd6544},
{-32'd1565, -32'd4671, 32'd10204, 32'd3398},
{32'd9453, -32'd6325, 32'd5052, -32'd2658},
{-32'd7680, 32'd5111, 32'd7686, 32'd2973},
{32'd8940, 32'd3662, 32'd8656, -32'd1265},
{-32'd14833, -32'd3660, 32'd2433, -32'd8591},
{32'd5693, -32'd4259, 32'd7957, -32'd10399},
{32'd12363, -32'd2295, 32'd8872, 32'd3460},
{32'd6804, -32'd5736, -32'd11872, 32'd2611},
{-32'd3796, 32'd11098, -32'd3475, -32'd5511},
{32'd776, 32'd9685, 32'd7444, -32'd5615},
{32'd111, -32'd4280, -32'd1452, -32'd711},
{-32'd8803, -32'd8968, -32'd6469, -32'd3935},
{-32'd2028, -32'd1613, -32'd6581, -32'd7269},
{-32'd9111, -32'd2592, 32'd5136, 32'd435},
{32'd5813, 32'd6805, 32'd4146, 32'd5510},
{32'd3124, 32'd1252, 32'd6873, 32'd1353},
{32'd1001, 32'd3006, 32'd5970, -32'd940},
{32'd1450, -32'd164, -32'd3071, -32'd2685},
{-32'd1003, -32'd9437, -32'd11179, 32'd10360},
{32'd1328, 32'd15705, -32'd3117, -32'd1072},
{-32'd8705, -32'd9308, 32'd1120, -32'd7487},
{-32'd268, 32'd7118, 32'd5434, -32'd1375},
{-32'd8002, -32'd5914, 32'd4291, 32'd4387},
{32'd10524, 32'd4210, -32'd6157, 32'd6319},
{-32'd4518, -32'd18541, -32'd12833, -32'd5812},
{32'd10493, -32'd5739, 32'd1168, 32'd4968},
{-32'd1408, 32'd10965, -32'd1481, -32'd8543},
{32'd3870, -32'd815, -32'd1735, -32'd4894},
{-32'd4282, 32'd3576, 32'd4187, 32'd2370},
{32'd8219, 32'd2949, -32'd492, -32'd2942},
{32'd914, 32'd5628, 32'd6378, 32'd5076},
{-32'd7487, 32'd7248, -32'd8557, -32'd3422},
{-32'd7151, -32'd3958, 32'd8169, 32'd7614},
{32'd6802, 32'd6981, 32'd2351, -32'd1910},
{-32'd1358, 32'd2431, 32'd1976, 32'd4039},
{32'd5994, -32'd8848, 32'd12454, 32'd4657},
{32'd6239, 32'd3591, -32'd2403, 32'd2063},
{-32'd8232, 32'd1653, -32'd8050, -32'd8506},
{-32'd5710, -32'd1281, -32'd3711, -32'd5362},
{32'd10951, -32'd814, -32'd6580, -32'd5355},
{-32'd1894, 32'd6722, -32'd7812, 32'd632},
{32'd1279, 32'd7245, 32'd3207, -32'd8190},
{-32'd1297, -32'd2215, -32'd3865, -32'd7726},
{-32'd3743, -32'd9200, 32'd2135, 32'd3977},
{32'd10061, -32'd5976, 32'd7095, 32'd5673},
{32'd6117, -32'd2213, -32'd5507, -32'd6388},
{32'd6471, -32'd125, 32'd1996, 32'd10009},
{-32'd6572, -32'd3695, 32'd4725, 32'd902},
{32'd13214, -32'd4518, -32'd9240, -32'd2214},
{-32'd2014, 32'd2076, -32'd3778, -32'd1977},
{-32'd16500, -32'd4081, -32'd1548, -32'd2177},
{32'd16604, -32'd407, 32'd11095, 32'd1232},
{32'd7312, 32'd2809, -32'd4380, 32'd317},
{32'd10743, 32'd1285, 32'd540, 32'd218},
{-32'd3632, 32'd12958, -32'd6797, -32'd2451},
{-32'd1255, -32'd10616, 32'd6904, 32'd4844},
{32'd1163, 32'd66, 32'd12298, -32'd3447},
{-32'd4119, 32'd7272, -32'd2836, -32'd2415},
{32'd1264, -32'd2882, -32'd10161, -32'd3944},
{32'd3777, 32'd6097, -32'd3421, -32'd2585},
{32'd11582, 32'd2072, 32'd9183, 32'd5285},
{32'd15293, -32'd7051, 32'd2190, -32'd143},
{-32'd249, -32'd2058, -32'd4352, -32'd1238},
{-32'd3076, -32'd1086, 32'd9121, -32'd4162},
{-32'd4487, -32'd2544, 32'd1491, 32'd2432},
{-32'd1441, -32'd7117, -32'd184, -32'd8464},
{-32'd2679, 32'd1184, 32'd8832, 32'd111},
{-32'd2418, -32'd8852, 32'd6853, 32'd2050},
{32'd6455, 32'd8568, 32'd3895, -32'd6604},
{-32'd7465, 32'd5934, -32'd210, -32'd743},
{-32'd3333, -32'd2013, -32'd9512, -32'd1074},
{32'd3230, -32'd743, -32'd867, -32'd207},
{-32'd5638, 32'd920, -32'd1303, -32'd6096},
{-32'd9779, -32'd5970, 32'd1455, -32'd6237},
{32'd8492, 32'd11187, -32'd791, -32'd5856},
{-32'd2296, 32'd2893, 32'd6886, 32'd4638},
{32'd547, 32'd1729, 32'd1732, 32'd1613},
{-32'd4843, -32'd2711, -32'd3878, -32'd5668},
{-32'd9905, 32'd2807, 32'd742, -32'd4736},
{32'd12205, -32'd2015, 32'd1091, 32'd8939},
{32'd1316, -32'd1087, -32'd5669, 32'd3667},
{32'd2662, -32'd17609, -32'd6035, 32'd527},
{-32'd7456, -32'd4715, 32'd5512, 32'd1794},
{32'd8031, 32'd5654, -32'd7859, -32'd3881},
{32'd4164, -32'd3615, -32'd2056, -32'd573},
{-32'd3903, -32'd3888, 32'd878, -32'd2490},
{32'd10744, 32'd2388, 32'd4168, -32'd2069},
{-32'd658, 32'd14302, -32'd3821, 32'd10072},
{-32'd4669, -32'd3306, -32'd9964, 32'd2297},
{-32'd9313, -32'd9585, -32'd3802, 32'd832},
{-32'd473, 32'd9653, 32'd4539, 32'd4482},
{-32'd4723, -32'd7219, 32'd6612, 32'd5555},
{-32'd3057, 32'd6362, 32'd840, -32'd8319},
{-32'd4950, -32'd14516, -32'd4896, -32'd1002},
{-32'd17357, 32'd2186, 32'd11497, -32'd5781},
{32'd5667, 32'd10350, 32'd11292, -32'd382},
{-32'd7089, 32'd2693, -32'd1454, 32'd4740},
{-32'd12403, -32'd884, -32'd5135, -32'd2704},
{32'd3116, -32'd12488, 32'd1068, 32'd2321},
{-32'd976, -32'd1084, 32'd5628, 32'd3178},
{-32'd9519, -32'd1414, -32'd5151, -32'd529},
{-32'd2328, -32'd7058, 32'd874, -32'd815},
{32'd5721, 32'd369, 32'd980, 32'd4271},
{-32'd1944, -32'd3668, -32'd1372, 32'd2717},
{32'd7612, 32'd8628, -32'd3271, -32'd14722},
{32'd6302, -32'd4679, -32'd3118, -32'd2029},
{-32'd4533, -32'd2707, -32'd8453, -32'd7514},
{-32'd1357, 32'd1566, 32'd6459, -32'd5013},
{-32'd8048, 32'd6362, -32'd5720, -32'd2318},
{-32'd4279, -32'd1811, 32'd5489, -32'd7049},
{-32'd7035, -32'd7200, 32'd5461, -32'd1769},
{32'd3010, 32'd5011, 32'd1992, -32'd2650},
{-32'd7887, 32'd2257, -32'd9462, -32'd8039},
{32'd751, -32'd2136, -32'd5315, -32'd5788},
{-32'd3125, -32'd1854, -32'd5703, -32'd1826},
{32'd7779, -32'd7595, 32'd10168, -32'd1178},
{-32'd5029, 32'd5657, -32'd6193, -32'd9087},
{-32'd6325, 32'd1717, 32'd4769, -32'd1671},
{32'd7257, -32'd743, 32'd3713, -32'd4756},
{-32'd5276, -32'd2850, 32'd1958, -32'd2443},
{-32'd8269, 32'd6650, -32'd3704, -32'd233},
{-32'd3675, 32'd1385, -32'd6988, -32'd258},
{32'd2362, 32'd3401, 32'd4, -32'd534},
{-32'd8330, 32'd907, 32'd2079, -32'd1049},
{-32'd6367, -32'd8114, 32'd851, 32'd6674},
{-32'd2047, 32'd820, 32'd828, 32'd1988},
{-32'd4968, -32'd1868, -32'd1636, 32'd2508},
{-32'd1130, -32'd1313, -32'd13305, -32'd701},
{32'd191, 32'd4631, 32'd6676, 32'd15553},
{-32'd3357, -32'd5851, 32'd4958, 32'd4836},
{-32'd4206, -32'd1682, -32'd6261, 32'd4902},
{-32'd1055, -32'd8562, -32'd2215, -32'd2834},
{-32'd4896, -32'd5247, -32'd5342, -32'd1721},
{-32'd599, 32'd9511, 32'd1774, 32'd9195},
{32'd3802, 32'd2182, 32'd8605, 32'd5116},
{32'd1243, -32'd5374, 32'd3049, 32'd3175},
{-32'd9446, 32'd8816, -32'd8743, -32'd425},
{-32'd3642, 32'd8524, -32'd801, -32'd1302},
{-32'd5021, -32'd2793, 32'd10778, 32'd7676},
{32'd3041, -32'd11531, 32'd6264, 32'd917},
{-32'd449, -32'd2991, 32'd5118, 32'd3709},
{-32'd3589, -32'd5467, 32'd5155, 32'd6391},
{32'd3969, 32'd2867, 32'd9616, 32'd475},
{-32'd901, 32'd7627, -32'd1915, -32'd9690},
{32'd7516, -32'd2863, 32'd6118, 32'd5142},
{-32'd5479, 32'd5386, -32'd13075, -32'd3701},
{32'd4345, 32'd4253, -32'd1212, 32'd7092},
{32'd7138, -32'd9331, -32'd2609, -32'd58},
{-32'd397, -32'd6770, -32'd2684, 32'd1666},
{32'd8832, -32'd5550, -32'd2279, 32'd2415},
{32'd1196, -32'd6612, 32'd304, -32'd1328},
{-32'd9798, 32'd5376, 32'd3007, -32'd10704},
{-32'd18254, -32'd2514, -32'd4328, -32'd4087},
{-32'd3018, 32'd15474, -32'd4798, -32'd8609},
{-32'd12494, 32'd3417, -32'd8346, -32'd241},
{32'd4891, -32'd7165, 32'd4817, -32'd3658},
{32'd2426, 32'd5968, 32'd13273, 32'd4183},
{-32'd2949, 32'd3821, -32'd14974, 32'd715}
},
{{32'd10361, 32'd45, 32'd4381, 32'd9242},
{-32'd1455, -32'd4047, -32'd6303, -32'd5251},
{-32'd4335, 32'd4595, 32'd4848, 32'd1283},
{32'd3716, -32'd9605, -32'd4273, 32'd9039},
{32'd2989, -32'd11932, 32'd7633, -32'd797},
{-32'd15293, 32'd808, 32'd7978, 32'd15582},
{-32'd915, -32'd2109, -32'd1339, 32'd7407},
{32'd8967, -32'd4605, -32'd4236, -32'd8512},
{-32'd229, 32'd3236, 32'd623, 32'd1155},
{32'd8398, 32'd3858, 32'd7972, 32'd3258},
{32'd5924, -32'd1293, 32'd5539, 32'd9921},
{-32'd7751, 32'd439, 32'd9226, 32'd3866},
{32'd7525, 32'd2120, 32'd2171, 32'd3666},
{-32'd7572, -32'd9003, 32'd3998, -32'd9958},
{-32'd6892, -32'd7828, -32'd16017, -32'd4735},
{32'd2907, 32'd552, -32'd5018, 32'd566},
{32'd10296, 32'd3796, 32'd4879, 32'd3419},
{32'd4990, 32'd4826, -32'd179, -32'd1424},
{-32'd13428, 32'd4537, -32'd3690, 32'd403},
{-32'd643, -32'd1683, 32'd2096, 32'd2356},
{-32'd7579, 32'd848, 32'd1809, 32'd10576},
{-32'd7643, -32'd8950, -32'd4557, -32'd10918},
{32'd8271, -32'd8085, 32'd574, 32'd4389},
{-32'd6344, 32'd3839, -32'd7264, -32'd5592},
{32'd1578, 32'd2616, 32'd4361, 32'd1223},
{32'd1458, -32'd858, 32'd1421, 32'd3826},
{32'd10318, 32'd2010, 32'd537, -32'd2380},
{32'd6908, 32'd11483, 32'd1434, -32'd7464},
{32'd7518, -32'd7783, 32'd16372, 32'd7850},
{32'd6597, 32'd7685, -32'd1063, -32'd12913},
{-32'd2862, 32'd832, 32'd3606, 32'd3380},
{-32'd3634, -32'd5868, -32'd5956, -32'd3505},
{32'd5669, 32'd3699, 32'd6633, -32'd4674},
{32'd6288, 32'd1408, -32'd52, -32'd6434},
{32'd5496, 32'd4910, 32'd7161, -32'd635},
{-32'd5556, 32'd1063, 32'd6202, 32'd8019},
{-32'd3704, 32'd9466, 32'd16, -32'd861},
{-32'd7647, 32'd2547, -32'd1650, -32'd9991},
{32'd1344, 32'd8677, 32'd3531, -32'd6219},
{32'd10644, 32'd5908, 32'd6313, -32'd14588},
{-32'd8084, -32'd1298, -32'd8003, 32'd3748},
{32'd8768, 32'd410, 32'd10044, 32'd1059},
{32'd9627, 32'd11442, -32'd712, -32'd1913},
{-32'd2914, 32'd6521, -32'd12459, -32'd4315},
{-32'd1174, -32'd9307, -32'd2747, -32'd18371},
{-32'd6017, 32'd6704, 32'd3516, -32'd7326},
{-32'd2979, -32'd6457, -32'd3170, -32'd4724},
{32'd1290, -32'd10756, -32'd2311, -32'd8261},
{32'd977, -32'd1425, 32'd4433, 32'd7974},
{-32'd8939, -32'd7665, -32'd513, 32'd5962},
{32'd3042, 32'd2203, -32'd718, -32'd7279},
{-32'd3918, 32'd6075, -32'd3983, -32'd3991},
{-32'd1780, -32'd8096, -32'd5171, -32'd1625},
{32'd3244, -32'd9336, -32'd3509, 32'd7840},
{-32'd7076, 32'd3580, 32'd2599, -32'd4595},
{32'd4351, -32'd3594, -32'd1028, -32'd10},
{-32'd4005, 32'd3083, 32'd8466, -32'd3163},
{-32'd13126, -32'd5808, -32'd6643, -32'd1094},
{-32'd16228, -32'd3642, -32'd5352, -32'd2242},
{32'd5208, 32'd9288, 32'd4514, 32'd8630},
{-32'd6703, -32'd10729, 32'd879, 32'd9332},
{32'd6427, -32'd2940, -32'd3850, 32'd1260},
{-32'd4915, -32'd7142, -32'd4976, -32'd3570},
{-32'd4137, 32'd198, -32'd3318, 32'd10442},
{32'd11347, 32'd9249, -32'd2970, -32'd5998},
{32'd1787, 32'd3385, 32'd9218, -32'd3165},
{32'd2897, 32'd5533, -32'd10688, -32'd3103},
{32'd2003, -32'd13200, -32'd1229, -32'd5568},
{32'd6275, -32'd406, -32'd13618, -32'd6501},
{-32'd5957, 32'd2437, -32'd152, 32'd1322},
{-32'd1874, 32'd12217, 32'd2280, -32'd15065},
{32'd2650, 32'd11334, 32'd7262, -32'd10538},
{-32'd545, 32'd5185, -32'd4086, 32'd4208},
{32'd6011, 32'd6260, -32'd1028, 32'd9046},
{32'd7755, 32'd2156, 32'd8622, 32'd6354},
{-32'd1484, 32'd591, -32'd7028, -32'd7673},
{32'd147, 32'd2493, -32'd5709, -32'd5613},
{32'd4267, -32'd14873, -32'd12376, 32'd13315},
{32'd7093, 32'd3251, 32'd1075, -32'd8446},
{32'd6809, 32'd1109, 32'd5659, 32'd2569},
{-32'd4468, -32'd14818, 32'd3396, 32'd1852},
{32'd184, 32'd4634, 32'd9566, 32'd4604},
{-32'd1722, 32'd8916, 32'd221, 32'd4903},
{-32'd6452, 32'd4137, 32'd3470, 32'd7927},
{-32'd5439, -32'd6367, 32'd952, -32'd6889},
{32'd1767, 32'd1741, 32'd7565, -32'd11016},
{32'd3364, -32'd1642, 32'd7979, -32'd8909},
{-32'd10854, 32'd3961, -32'd1678, 32'd2707},
{-32'd4595, -32'd7257, -32'd9471, -32'd5295},
{32'd450, -32'd6712, -32'd5954, -32'd3978},
{32'd5736, 32'd1121, 32'd4420, 32'd113},
{32'd1057, 32'd683, -32'd3102, 32'd2802},
{32'd14241, -32'd5373, 32'd141, -32'd10151},
{-32'd2681, -32'd4435, 32'd5227, -32'd1074},
{32'd2404, 32'd397, -32'd8350, -32'd8922},
{-32'd4883, -32'd1679, -32'd1219, -32'd9435},
{-32'd3566, 32'd242, -32'd21, -32'd245},
{32'd4938, -32'd1318, 32'd1124, 32'd11176},
{-32'd7511, 32'd4301, 32'd2071, -32'd46},
{32'd13965, -32'd4577, 32'd13590, 32'd1524},
{-32'd82, -32'd1205, -32'd12205, 32'd5376},
{32'd861, 32'd1360, 32'd4488, -32'd4519},
{32'd642, 32'd3955, -32'd6585, -32'd374},
{32'd11065, 32'd5021, -32'd693, 32'd10802},
{32'd3885, 32'd15340, 32'd6144, 32'd632},
{-32'd1658, -32'd12126, 32'd5019, 32'd7830},
{32'd1416, -32'd1985, -32'd249, 32'd3756},
{32'd7625, -32'd6011, 32'd3520, -32'd436},
{32'd9507, 32'd3326, 32'd2797, 32'd9935},
{-32'd397, 32'd1007, -32'd703, 32'd254},
{-32'd6426, -32'd5197, -32'd9772, 32'd367},
{32'd3728, 32'd7738, -32'd1928, -32'd5461},
{32'd14099, -32'd645, -32'd346, 32'd10194},
{-32'd8567, 32'd2954, 32'd7526, 32'd1901},
{-32'd7261, -32'd11097, -32'd5850, 32'd1102},
{-32'd5566, -32'd9627, 32'd1378, 32'd7643},
{32'd6948, 32'd2591, 32'd10691, 32'd4836},
{32'd11557, -32'd5188, 32'd1843, -32'd14510},
{32'd4847, -32'd1468, 32'd6060, -32'd1552},
{32'd6930, -32'd3545, 32'd6800, 32'd6269},
{32'd4096, 32'd3820, -32'd3739, -32'd5355},
{-32'd1769, -32'd2388, -32'd4599, 32'd4600},
{-32'd2771, 32'd2112, 32'd1433, -32'd11196},
{-32'd5925, -32'd5644, 32'd9540, -32'd5719},
{32'd2480, 32'd7140, -32'd1109, 32'd3730},
{32'd3190, -32'd499, 32'd8452, 32'd4261},
{32'd1598, -32'd12614, 32'd5, 32'd7875},
{32'd1199, 32'd3280, -32'd4463, -32'd8012},
{32'd2638, 32'd4860, -32'd5947, 32'd3725},
{-32'd7727, 32'd1980, -32'd477, 32'd2041},
{-32'd6239, -32'd116, -32'd723, 32'd6950},
{-32'd5672, -32'd537, -32'd517, -32'd3725},
{-32'd5192, 32'd2197, -32'd10724, 32'd2445},
{-32'd3375, 32'd9605, -32'd879, -32'd7159},
{32'd4027, 32'd7379, 32'd4936, -32'd5477},
{32'd11804, 32'd1681, 32'd8943, -32'd5313},
{-32'd4428, -32'd6897, -32'd1964, -32'd8564},
{-32'd552, -32'd1931, -32'd9278, 32'd1594},
{32'd2968, -32'd4610, 32'd3460, -32'd1918},
{-32'd4663, -32'd3932, -32'd5339, -32'd3464},
{32'd112, 32'd1741, -32'd8264, 32'd5529},
{-32'd7556, -32'd3941, 32'd482, -32'd15345},
{32'd3905, -32'd4745, 32'd7702, 32'd2802},
{32'd7291, 32'd3107, 32'd2180, 32'd7808},
{32'd1291, 32'd11630, 32'd9962, -32'd1280},
{-32'd4628, 32'd6130, -32'd5693, -32'd6616},
{-32'd4695, -32'd622, 32'd12555, -32'd5024},
{32'd838, 32'd7656, 32'd7211, -32'd9473},
{32'd1006, 32'd2443, 32'd3965, -32'd625},
{-32'd11207, -32'd6616, -32'd5770, -32'd2969},
{32'd636, 32'd520, -32'd4782, -32'd4468},
{-32'd4103, -32'd6549, 32'd3142, 32'd6311},
{-32'd6816, -32'd5984, 32'd1208, -32'd1277},
{-32'd245, 32'd6618, 32'd4605, 32'd258},
{32'd292, 32'd4187, 32'd533, -32'd13619},
{32'd6283, 32'd329, -32'd7081, -32'd12774},
{32'd1556, 32'd3210, 32'd9542, 32'd9222},
{-32'd2817, 32'd5787, 32'd6253, 32'd4958},
{-32'd4347, -32'd14687, -32'd9073, 32'd7160},
{-32'd5, -32'd6515, -32'd267, -32'd6064},
{-32'd11879, -32'd4051, -32'd28, 32'd3251},
{-32'd211, -32'd6374, 32'd3231, 32'd3018},
{32'd4398, -32'd2478, 32'd3988, 32'd1313},
{-32'd4350, 32'd7042, 32'd4116, 32'd688},
{32'd699, 32'd10907, 32'd3698, -32'd592},
{-32'd3697, 32'd12026, -32'd8618, 32'd1355},
{32'd3680, 32'd1479, -32'd1694, -32'd2519},
{-32'd12221, 32'd1089, 32'd500, -32'd7179},
{-32'd8077, 32'd1236, -32'd15, -32'd5174},
{-32'd608, 32'd6659, -32'd1028, -32'd2761},
{-32'd4069, -32'd3036, 32'd172, -32'd357},
{-32'd2177, 32'd4365, -32'd3013, 32'd1480},
{32'd13179, 32'd4392, 32'd6811, 32'd1884},
{-32'd7458, -32'd11500, -32'd4640, -32'd9006},
{32'd4047, -32'd3194, 32'd6872, -32'd171},
{32'd7655, 32'd9715, -32'd1538, -32'd4475},
{32'd8852, 32'd102, 32'd7357, 32'd6949},
{-32'd5071, 32'd601, -32'd3408, -32'd2970},
{32'd5068, -32'd1200, 32'd8113, 32'd5384},
{-32'd6031, -32'd4303, -32'd9254, -32'd6181},
{-32'd1057, -32'd3974, -32'd2344, 32'd2621},
{-32'd5796, -32'd10016, 32'd12403, 32'd2509},
{-32'd8501, 32'd4845, -32'd9043, -32'd3801},
{32'd1382, 32'd5069, -32'd1793, -32'd11935},
{32'd1432, -32'd12, 32'd7286, -32'd4671},
{32'd565, -32'd5523, 32'd4496, 32'd11382},
{-32'd58, 32'd594, 32'd6153, -32'd4500},
{32'd7406, -32'd1920, 32'd11966, 32'd7859},
{-32'd6968, 32'd2641, -32'd981, 32'd3084},
{-32'd7802, -32'd190, -32'd1616, 32'd2397},
{32'd5798, -32'd1111, -32'd11133, -32'd7367},
{-32'd6617, 32'd1399, -32'd9376, -32'd4835},
{-32'd5972, -32'd8089, -32'd3486, -32'd691},
{32'd1114, 32'd2263, -32'd1510, -32'd1669},
{32'd1522, -32'd7713, 32'd5585, 32'd3478},
{32'd2713, -32'd5679, 32'd5991, 32'd9568},
{32'd2512, 32'd3710, 32'd4701, 32'd12189},
{32'd11092, 32'd14724, 32'd11878, -32'd4807},
{-32'd3043, -32'd12775, 32'd14036, -32'd3800},
{-32'd6470, -32'd1803, -32'd938, -32'd6869},
{-32'd9560, -32'd6242, -32'd9003, -32'd3235},
{32'd869, 32'd3381, -32'd11486, -32'd4436},
{-32'd15297, 32'd5912, 32'd10524, 32'd340},
{-32'd4997, -32'd3886, 32'd2334, 32'd2084},
{-32'd11982, 32'd5815, -32'd7526, 32'd3544},
{-32'd1090, 32'd5188, 32'd2727, -32'd4785},
{32'd11548, 32'd94, 32'd8348, 32'd10376},
{-32'd1063, 32'd1429, -32'd8908, -32'd8316},
{-32'd3507, -32'd5184, -32'd3172, -32'd7611},
{32'd2296, 32'd8012, -32'd2345, -32'd21140},
{-32'd1062, 32'd3466, -32'd1276, -32'd9260},
{-32'd6720, -32'd910, -32'd3900, -32'd1231},
{32'd745, -32'd4450, 32'd5312, -32'd8675},
{32'd6373, -32'd2602, -32'd13177, 32'd1068},
{-32'd13328, 32'd2120, -32'd414, -32'd15533},
{-32'd9227, -32'd2890, -32'd5673, 32'd1079},
{32'd3267, 32'd6719, 32'd3522, -32'd10151},
{-32'd2989, 32'd3783, -32'd3601, -32'd14502},
{-32'd2519, 32'd11510, 32'd5295, -32'd5704},
{32'd2358, 32'd703, -32'd8778, -32'd8942},
{32'd8731, -32'd4166, -32'd836, 32'd2389},
{-32'd1107, -32'd3350, -32'd1165, 32'd12147},
{32'd2738, -32'd15383, 32'd1280, 32'd8735},
{-32'd657, 32'd5895, 32'd4732, 32'd6},
{-32'd269, 32'd749, 32'd3822, 32'd13599},
{-32'd8515, 32'd401, 32'd1683, 32'd2938},
{32'd10096, -32'd5002, -32'd10700, 32'd5617},
{-32'd11189, -32'd3747, 32'd607, 32'd6262},
{-32'd1229, -32'd2482, -32'd991, -32'd4239},
{32'd105, 32'd2662, 32'd4323, 32'd589},
{32'd8744, -32'd1451, -32'd3235, -32'd13389},
{32'd10509, -32'd6011, 32'd4193, 32'd2574},
{-32'd3841, -32'd5197, -32'd281, 32'd18439},
{32'd5207, -32'd1370, 32'd8647, 32'd615},
{32'd4794, 32'd1640, -32'd6096, -32'd5974},
{-32'd6254, 32'd3018, -32'd8445, -32'd9810},
{32'd7140, -32'd7304, 32'd12461, -32'd6597},
{32'd4739, 32'd2841, -32'd2975, 32'd573},
{-32'd1168, 32'd3661, -32'd3015, 32'd9276},
{-32'd11708, 32'd9733, -32'd4823, -32'd1895},
{32'd3504, 32'd3881, 32'd1696, -32'd1036},
{32'd14184, 32'd1674, 32'd688, -32'd6440},
{32'd1854, -32'd1114, -32'd3569, -32'd7310},
{-32'd2299, 32'd7707, -32'd873, -32'd3690},
{32'd16909, 32'd2985, 32'd5294, 32'd12496},
{-32'd11115, -32'd4333, -32'd7986, 32'd7679},
{-32'd8047, 32'd5015, -32'd4988, -32'd16552},
{32'd4069, -32'd2262, 32'd8417, -32'd3766},
{-32'd1317, 32'd4255, 32'd1876, -32'd780},
{32'd5570, 32'd10434, 32'd4841, -32'd4622},
{32'd311, -32'd182, 32'd1723, 32'd6625},
{32'd1402, 32'd1179, -32'd5102, -32'd8455},
{32'd2687, -32'd7564, -32'd3717, -32'd6546},
{-32'd3487, 32'd6594, -32'd12441, 32'd2331},
{-32'd11499, -32'd5964, -32'd9257, 32'd2308},
{-32'd6114, 32'd5711, 32'd7346, -32'd4382},
{-32'd203, -32'd5177, -32'd2543, 32'd7027},
{32'd7166, 32'd6240, -32'd8540, -32'd5259},
{-32'd10457, 32'd7881, -32'd4653, -32'd1472},
{32'd541, 32'd8047, 32'd187, -32'd5777},
{32'd8087, -32'd6163, 32'd684, 32'd2926},
{32'd699, 32'd4748, -32'd6833, 32'd7627},
{-32'd13079, -32'd18891, -32'd7751, 32'd2829},
{32'd5171, -32'd3950, -32'd7785, -32'd5177},
{32'd4814, -32'd3094, 32'd679, 32'd8779},
{-32'd2162, 32'd4668, 32'd5205, 32'd1175},
{32'd8421, -32'd4222, 32'd409, 32'd12094},
{-32'd920, 32'd9288, 32'd4708, 32'd8371},
{-32'd13611, -32'd2039, -32'd162, 32'd3460},
{32'd10, -32'd5364, -32'd1999, -32'd46},
{32'd4017, 32'd2837, -32'd5081, 32'd7327},
{-32'd1869, 32'd4979, 32'd7032, 32'd11553},
{-32'd6297, -32'd3560, -32'd248, 32'd6228},
{-32'd5160, -32'd46, 32'd899, 32'd4015},
{-32'd7038, -32'd5951, -32'd432, 32'd3199},
{-32'd4813, -32'd63, 32'd3567, 32'd4929},
{32'd12466, 32'd5203, 32'd10496, 32'd4963},
{32'd1434, -32'd703, -32'd6155, -32'd3009},
{-32'd10898, -32'd5838, -32'd6584, 32'd3692},
{32'd6082, 32'd5324, -32'd3658, -32'd2910},
{32'd8107, -32'd2098, 32'd3033, -32'd2142},
{32'd19456, 32'd12370, 32'd9541, -32'd6059},
{32'd6824, -32'd4068, 32'd1678, 32'd5868},
{32'd1623, 32'd6722, -32'd211, -32'd2401},
{32'd7583, 32'd4888, 32'd17524, 32'd5236},
{-32'd14319, -32'd3760, -32'd8095, 32'd52},
{32'd601, 32'd3539, 32'd2332, 32'd10824},
{-32'd1694, -32'd4208, -32'd2631, 32'd2121},
{-32'd91, -32'd2038, 32'd2667, -32'd7182},
{32'd6273, -32'd3580, -32'd4535, 32'd8261},
{-32'd1428, -32'd5507, 32'd4047, 32'd10095},
{32'd6270, 32'd8246, 32'd11223, 32'd16541},
{-32'd1773, 32'd839, -32'd291, 32'd8377},
{-32'd4602, -32'd3793, -32'd1249, 32'd5210},
{-32'd7552, 32'd7591, -32'd5582, -32'd22},
{-32'd483, 32'd1312, -32'd2637, -32'd17822},
{-32'd8424, -32'd6847, -32'd2628, 32'd8265},
{32'd13073, -32'd6696, 32'd3905, -32'd5316},
{32'd976, 32'd1239, -32'd122, -32'd10137},
{-32'd13533, 32'd5766, -32'd6519, 32'd12474}
},
{{-32'd11775, -32'd931, -32'd1564, -32'd1825},
{32'd1353, 32'd2465, 32'd9451, -32'd4349},
{32'd5768, -32'd439, 32'd2027, -32'd9692},
{32'd7343, 32'd9844, -32'd4699, 32'd14500},
{32'd871, -32'd15431, -32'd2920, 32'd10834},
{32'd1427, 32'd5003, -32'd1299, 32'd5724},
{32'd9225, 32'd5200, -32'd3329, 32'd15215},
{32'd6295, -32'd8374, 32'd7713, -32'd9692},
{-32'd6667, -32'd3958, 32'd25447, -32'd4293},
{-32'd1572, 32'd5100, -32'd3385, 32'd13564},
{32'd12048, -32'd7374, -32'd1616, 32'd4921},
{-32'd7550, 32'd3882, 32'd1022, -32'd2907},
{-32'd1202, 32'd6695, -32'd6885, -32'd7338},
{-32'd5297, 32'd304, 32'd4674, 32'd9204},
{-32'd4934, 32'd12014, -32'd3288, -32'd12244},
{-32'd16684, -32'd8639, 32'd11810, 32'd60},
{32'd5197, 32'd2288, 32'd2051, -32'd8079},
{-32'd7523, 32'd7688, -32'd30, -32'd5032},
{-32'd466, -32'd3925, -32'd14759, 32'd2300},
{-32'd4914, 32'd3855, -32'd4, 32'd6111},
{-32'd6866, 32'd2455, -32'd9062, -32'd6408},
{-32'd11851, 32'd2943, -32'd9936, 32'd5124},
{32'd4828, 32'd1505, 32'd11270, -32'd10993},
{-32'd2136, 32'd3823, -32'd11447, -32'd2862},
{-32'd4814, 32'd5062, -32'd9226, 32'd5271},
{32'd1545, -32'd2681, -32'd271, 32'd291},
{32'd7987, -32'd8730, -32'd8840, 32'd201},
{32'd14064, 32'd4457, 32'd4439, 32'd503},
{32'd11411, 32'd5387, 32'd13957, 32'd8115},
{-32'd8188, -32'd13444, -32'd2969, -32'd191},
{-32'd2420, -32'd5182, -32'd7988, 32'd9919},
{-32'd7603, 32'd4496, -32'd9937, 32'd4541},
{-32'd3348, -32'd4680, -32'd3881, 32'd5164},
{32'd4871, -32'd11055, 32'd3270, 32'd521},
{32'd2284, 32'd8151, -32'd6564, 32'd4135},
{-32'd11328, -32'd8052, -32'd4045, -32'd3232},
{32'd8405, -32'd685, -32'd1357, -32'd2157},
{-32'd1036, -32'd5202, 32'd11054, 32'd448},
{32'd18957, 32'd14283, -32'd5981, 32'd2022},
{32'd3912, 32'd5244, 32'd2071, 32'd4008},
{32'd1794, 32'd10585, -32'd712, -32'd5162},
{-32'd2182, -32'd2968, -32'd6388, -32'd4651},
{-32'd3771, -32'd2987, -32'd3786, 32'd5871},
{-32'd1684, -32'd5534, -32'd1618, -32'd2085},
{-32'd24438, -32'd1506, 32'd5560, -32'd3753},
{-32'd10705, 32'd11473, -32'd40, 32'd7899},
{-32'd621, 32'd692, -32'd9764, -32'd4895},
{-32'd2076, -32'd7137, -32'd3419, 32'd2507},
{32'd6670, -32'd2710, -32'd2967, -32'd6724},
{-32'd9826, -32'd4356, 32'd745, -32'd5625},
{-32'd2728, -32'd10962, 32'd12540, -32'd1311},
{-32'd5266, 32'd12900, -32'd8106, -32'd1185},
{-32'd4285, 32'd4504, 32'd1284, -32'd3837},
{-32'd4349, -32'd2429, -32'd5268, -32'd12437},
{-32'd6586, -32'd11637, 32'd4129, 32'd1732},
{32'd8035, 32'd2091, 32'd18129, 32'd2662},
{32'd19945, 32'd2302, -32'd4763, 32'd1433},
{-32'd7201, -32'd4238, 32'd5883, 32'd2492},
{-32'd7919, 32'd3324, -32'd3378, -32'd2748},
{-32'd7962, 32'd2045, -32'd5496, 32'd987},
{32'd8250, 32'd2661, 32'd9096, -32'd3895},
{32'd13309, -32'd4891, -32'd6353, -32'd3991},
{-32'd8743, -32'd6118, 32'd9338, -32'd3727},
{-32'd8533, 32'd1904, -32'd10044, 32'd9577},
{-32'd3009, -32'd4829, -32'd3693, -32'd960},
{32'd8519, 32'd3300, -32'd4883, -32'd3814},
{32'd4042, 32'd3281, 32'd14169, 32'd2683},
{32'd13431, 32'd325, 32'd11838, -32'd9210},
{-32'd12206, 32'd1694, -32'd8154, 32'd3341},
{32'd10458, 32'd2276, 32'd5815, -32'd1997},
{-32'd640, 32'd1514, 32'd10377, 32'd5028},
{32'd20351, 32'd5168, 32'd7798, -32'd720},
{-32'd13437, -32'd2454, -32'd7863, -32'd8747},
{32'd14068, -32'd4733, 32'd8160, -32'd5943},
{32'd8378, 32'd4791, 32'd2370, -32'd321},
{32'd3089, 32'd789, -32'd3495, -32'd14263},
{32'd4143, -32'd5464, 32'd4369, -32'd5103},
{-32'd1171, -32'd7527, -32'd6336, -32'd5534},
{32'd7302, -32'd809, -32'd6406, -32'd3899},
{32'd5296, 32'd259, 32'd12008, 32'd10838},
{32'd3222, -32'd5027, -32'd9190, -32'd1097},
{-32'd4275, 32'd38, -32'd15750, 32'd3088},
{32'd3450, -32'd981, 32'd6322, 32'd6993},
{32'd5364, 32'd385, 32'd10676, 32'd840},
{-32'd9237, -32'd3345, 32'd2199, -32'd1681},
{32'd8659, -32'd2375, 32'd5077, 32'd10965},
{-32'd8839, 32'd19, -32'd11335, 32'd342},
{-32'd3736, -32'd1422, 32'd4098, 32'd8629},
{32'd7117, -32'd3177, 32'd11090, -32'd2063},
{-32'd10453, 32'd2219, 32'd10741, 32'd3910},
{32'd1097, 32'd7050, 32'd2468, 32'd1695},
{32'd10651, -32'd1695, -32'd5187, -32'd7946},
{32'd5733, -32'd1105, -32'd7693, 32'd9021},
{32'd12474, 32'd134, 32'd717, 32'd5227},
{32'd8520, -32'd6068, -32'd568, 32'd3045},
{-32'd7244, 32'd49, 32'd6076, 32'd8946},
{-32'd818, 32'd359, -32'd14141, 32'd7641},
{-32'd16102, -32'd4897, 32'd19603, -32'd4178},
{32'd3616, 32'd11696, 32'd1426, 32'd4929},
{-32'd7120, 32'd2701, -32'd4594, 32'd8172},
{-32'd2041, -32'd7019, -32'd628, 32'd2920},
{32'd4908, 32'd4690, -32'd2803, -32'd5117},
{-32'd1553, 32'd4894, 32'd3238, 32'd9812},
{-32'd32, -32'd1186, 32'd440, -32'd4298},
{32'd18897, -32'd1035, -32'd2762, 32'd4540},
{-32'd8275, -32'd10684, -32'd10630, -32'd542},
{-32'd914, 32'd8667, 32'd2, -32'd5959},
{-32'd931, -32'd7699, 32'd14490, -32'd8096},
{-32'd3007, -32'd3775, -32'd17103, -32'd4063},
{-32'd2061, -32'd6682, 32'd11664, -32'd6009},
{-32'd3126, 32'd10183, 32'd359, -32'd1856},
{-32'd10261, 32'd1391, -32'd12875, 32'd4222},
{32'd9894, 32'd1129, -32'd9014, -32'd25},
{-32'd4012, -32'd1810, -32'd15282, -32'd7425},
{-32'd5104, -32'd1486, -32'd8399, -32'd3519},
{32'd7211, -32'd211, 32'd12030, -32'd14720},
{32'd7972, 32'd2542, -32'd10435, -32'd11587},
{-32'd3440, 32'd8810, 32'd3972, -32'd10893},
{-32'd4587, 32'd3810, 32'd9943, 32'd14034},
{-32'd2556, 32'd6304, -32'd2486, -32'd4076},
{32'd13226, 32'd820, -32'd8008, 32'd2057},
{32'd14338, -32'd3136, -32'd18318, 32'd5514},
{32'd5246, 32'd201, 32'd7162, -32'd7704},
{32'd2119, 32'd12706, 32'd17346, 32'd3871},
{-32'd16651, -32'd11324, -32'd14841, -32'd13145},
{32'd2269, -32'd4437, 32'd14085, -32'd4052},
{32'd2220, -32'd228, -32'd8905, -32'd4806},
{32'd335, 32'd3367, 32'd774, -32'd5220},
{32'd840, -32'd7552, 32'd6208, 32'd9343},
{-32'd2632, 32'd2849, 32'd178, -32'd6078},
{-32'd10696, 32'd12500, -32'd13258, 32'd5048},
{-32'd701, -32'd6381, 32'd12620, -32'd5689},
{-32'd3033, -32'd1721, -32'd885, 32'd6657},
{32'd10584, -32'd3260, 32'd4595, 32'd1953},
{-32'd4431, 32'd2147, 32'd2993, 32'd12387},
{-32'd5369, 32'd1004, 32'd5822, 32'd6885},
{32'd7315, 32'd6489, 32'd14484, 32'd12526},
{-32'd6561, 32'd9086, -32'd8637, 32'd6765},
{-32'd6156, 32'd1523, 32'd10329, -32'd4595},
{-32'd5966, -32'd7961, -32'd1056, -32'd1661},
{-32'd4578, -32'd12828, -32'd8173, 32'd2327},
{-32'd3505, 32'd6398, 32'd7474, -32'd1220},
{-32'd2047, 32'd4166, -32'd7431, -32'd9403},
{-32'd5473, -32'd3288, 32'd12919, 32'd9499},
{32'd10098, 32'd267, -32'd7636, 32'd6589},
{32'd14921, 32'd5962, 32'd6250, 32'd832},
{32'd4072, -32'd354, -32'd14358, 32'd4876},
{-32'd8184, 32'd9794, -32'd17693, -32'd5242},
{-32'd664, 32'd7049, 32'd7892, 32'd12525},
{-32'd7091, 32'd8726, -32'd7449, -32'd12860},
{-32'd533, -32'd5330, 32'd294, -32'd9706},
{-32'd3737, 32'd2508, 32'd7477, -32'd7148},
{-32'd13478, -32'd6569, 32'd1090, -32'd6843},
{32'd2516, -32'd4720, -32'd1545, -32'd3417},
{32'd2360, 32'd8249, 32'd1479, -32'd14485},
{-32'd2874, 32'd14191, -32'd1306, 32'd6633},
{32'd1649, -32'd9960, -32'd9229, 32'd7128},
{32'd7718, 32'd7898, -32'd5654, -32'd7479},
{32'd9749, 32'd5663, -32'd10093, 32'd36},
{-32'd20107, -32'd4916, -32'd6707, -32'd142},
{-32'd10335, -32'd3299, -32'd153, -32'd19262},
{-32'd2793, -32'd4141, 32'd5443, -32'd622},
{32'd489, 32'd242, -32'd13276, -32'd5124},
{-32'd5638, 32'd10501, 32'd8085, 32'd2179},
{-32'd390, -32'd2368, 32'd2827, 32'd7242},
{-32'd18421, 32'd23156, 32'd7952, 32'd1125},
{32'd3358, -32'd1168, 32'd3817, 32'd8870},
{-32'd1682, 32'd4001, 32'd2328, -32'd6373},
{-32'd3090, -32'd6776, -32'd9990, 32'd2720},
{32'd1704, -32'd8085, 32'd12064, -32'd4202},
{32'd10021, 32'd5613, 32'd403, 32'd9007},
{32'd5549, 32'd845, -32'd5654, 32'd4517},
{-32'd2825, 32'd10855, 32'd1842, 32'd8020},
{32'd6670, -32'd11960, -32'd6432, -32'd2403},
{32'd1697, -32'd4392, 32'd3788, -32'd4756},
{-32'd9748, -32'd9582, 32'd1941, -32'd1664},
{-32'd1359, -32'd4749, 32'd2513, 32'd4634},
{32'd9088, 32'd18340, 32'd10734, 32'd4240},
{-32'd1226, 32'd8343, 32'd795, 32'd5330},
{32'd1, -32'd4538, 32'd3761, -32'd13741},
{-32'd4862, 32'd6747, 32'd4445, 32'd1611},
{-32'd4357, -32'd11022, 32'd4662, 32'd1765},
{-32'd4320, 32'd3447, -32'd2298, -32'd1781},
{-32'd14841, -32'd7211, 32'd782, 32'd6384},
{32'd1229, -32'd13821, 32'd2652, 32'd7474},
{32'd4019, 32'd6932, 32'd5208, 32'd1400},
{-32'd1208, 32'd17133, 32'd3639, -32'd6731},
{32'd7787, 32'd147, 32'd5759, -32'd9590},
{32'd10168, -32'd3106, 32'd13795, 32'd5041},
{-32'd11023, 32'd201, 32'd948, 32'd2569},
{-32'd379, -32'd4021, -32'd7552, 32'd2638},
{32'd4069, -32'd147, 32'd981, -32'd1274},
{32'd5073, -32'd3842, 32'd5927, 32'd16236},
{-32'd1280, -32'd2987, -32'd19728, -32'd8774},
{-32'd2636, -32'd1154, 32'd17742, -32'd78},
{-32'd8619, 32'd77, -32'd12644, -32'd11332},
{-32'd9093, -32'd7776, 32'd3898, -32'd3556},
{32'd13236, -32'd4525, 32'd4279, -32'd1036},
{32'd4507, 32'd3616, 32'd6405, 32'd5013},
{-32'd10747, 32'd8504, -32'd8003, 32'd338},
{-32'd2731, -32'd2293, -32'd5256, -32'd4671},
{32'd3096, 32'd6447, -32'd5828, 32'd7943},
{32'd4492, -32'd1324, -32'd1902, 32'd8207},
{32'd28631, 32'd10747, 32'd6442, -32'd6955},
{32'd144, -32'd9076, 32'd3470, 32'd5598},
{32'd13505, 32'd14967, 32'd9393, -32'd3312},
{-32'd8349, -32'd4095, 32'd12393, 32'd7091},
{32'd16531, 32'd7157, 32'd4855, 32'd12701},
{32'd9730, -32'd5827, 32'd9492, 32'd4962},
{32'd8852, -32'd3544, -32'd3144, 32'd13327},
{32'd2018, -32'd6944, 32'd5783, -32'd19480},
{-32'd3833, 32'd3859, -32'd3900, 32'd4445},
{-32'd11518, -32'd2760, 32'd7130, 32'd4387},
{-32'd3872, -32'd2548, 32'd11331, 32'd6654},
{-32'd14513, -32'd1191, -32'd8834, -32'd6504},
{32'd5439, -32'd2686, -32'd3567, -32'd3121},
{32'd750, 32'd7861, 32'd19380, -32'd2845},
{-32'd1401, -32'd7265, 32'd8329, 32'd2242},
{32'd13513, 32'd7072, -32'd4070, 32'd10287},
{32'd361, 32'd12669, 32'd1797, -32'd4820},
{-32'd1859, 32'd4282, 32'd22692, -32'd2208},
{32'd2272, -32'd288, -32'd3734, 32'd11547},
{32'd921, 32'd107, -32'd1816, -32'd2496},
{-32'd12555, 32'd11202, -32'd2875, -32'd1046},
{-32'd3385, -32'd8858, -32'd5238, 32'd4647},
{-32'd2965, -32'd6252, 32'd3384, -32'd3942},
{32'd4357, -32'd426, 32'd12140, 32'd1892},
{-32'd2111, -32'd8635, -32'd1691, 32'd1041},
{32'd5725, 32'd6357, -32'd3952, -32'd2182},
{32'd12386, 32'd6216, -32'd2604, 32'd1070},
{-32'd7212, -32'd7570, -32'd9233, -32'd10808},
{32'd8932, -32'd383, 32'd864, -32'd112},
{-32'd576, 32'd2227, -32'd8204, 32'd866},
{-32'd217, -32'd7638, -32'd3387, -32'd7976},
{-32'd4729, 32'd1987, 32'd10149, -32'd6758},
{32'd9492, 32'd1398, 32'd9283, -32'd6719},
{32'd1733, 32'd8716, 32'd15564, 32'd532},
{32'd5680, -32'd10249, -32'd361, 32'd7293},
{32'd1122, 32'd3275, -32'd804, -32'd1541},
{-32'd1058, 32'd7048, 32'd9023, 32'd1083},
{32'd11505, -32'd1652, -32'd15925, -32'd937},
{-32'd8951, -32'd11938, 32'd5505, -32'd5357},
{32'd26, -32'd2794, 32'd1173, -32'd7177},
{32'd10585, -32'd5643, 32'd9181, 32'd1466},
{-32'd216, 32'd1226, -32'd1490, 32'd6866},
{-32'd2973, -32'd2488, -32'd18454, -32'd3610},
{32'd6015, -32'd4697, 32'd4759, 32'd6003},
{-32'd4948, -32'd719, -32'd1110, 32'd5505},
{-32'd490, -32'd6433, -32'd7366, -32'd6018},
{32'd10739, -32'd4048, -32'd4262, 32'd1615},
{-32'd981, -32'd13334, 32'd7002, 32'd6094},
{-32'd1704, 32'd4303, -32'd5307, -32'd7316},
{-32'd403, 32'd992, 32'd7202, 32'd4468},
{32'd2219, -32'd3144, -32'd5385, 32'd990},
{-32'd3927, -32'd492, 32'd10650, -32'd4806},
{32'd2854, 32'd11380, 32'd6256, 32'd1390},
{32'd4784, -32'd5235, -32'd7482, 32'd789},
{-32'd6420, 32'd5139, -32'd6693, 32'd7406},
{-32'd3020, -32'd3960, -32'd8364, -32'd400},
{-32'd2803, -32'd3417, 32'd10961, -32'd7348},
{32'd6928, 32'd1313, 32'd15700, -32'd4978},
{32'd1584, -32'd2214, 32'd554, -32'd6777},
{-32'd5753, -32'd5442, -32'd1322, -32'd3701},
{32'd5375, 32'd4459, -32'd6446, -32'd5063},
{32'd7020, 32'd5852, 32'd19830, -32'd6715},
{-32'd3149, 32'd12246, -32'd16069, -32'd2887},
{-32'd4308, 32'd9053, -32'd6810, 32'd7584},
{-32'd4119, -32'd3872, -32'd6733, -32'd8965},
{-32'd2574, -32'd2891, -32'd81, 32'd708},
{32'd8896, -32'd4227, 32'd3507, -32'd5365},
{-32'd2667, 32'd6795, 32'd11381, -32'd4224},
{32'd569, 32'd272, 32'd2219, -32'd2325},
{32'd6014, 32'd3864, -32'd97, -32'd4618},
{-32'd18252, 32'd2826, 32'd20379, -32'd8417},
{-32'd4225, -32'd1111, 32'd2598, -32'd5060},
{32'd11215, -32'd9769, -32'd1951, -32'd9986},
{32'd1084, 32'd6996, -32'd481, 32'd8754},
{32'd7299, 32'd8424, 32'd844, 32'd8211},
{-32'd5139, -32'd10010, 32'd4055, -32'd7130},
{32'd5335, -32'd6263, -32'd7119, 32'd1184},
{-32'd1146, 32'd8085, -32'd1632, 32'd10680},
{-32'd6940, -32'd4630, 32'd11515, -32'd1081},
{32'd5432, 32'd5186, 32'd13945, 32'd16415},
{32'd17590, -32'd3444, -32'd942, 32'd10974},
{-32'd2746, 32'd2416, 32'd4187, -32'd3924},
{-32'd5392, -32'd7198, 32'd1364, 32'd308},
{32'd246, 32'd5481, 32'd5473, 32'd6885},
{-32'd12199, -32'd4125, -32'd4205, -32'd6420},
{-32'd1787, -32'd395, 32'd1483, -32'd4225},
{32'd11509, 32'd6711, -32'd13767, -32'd9668},
{32'd3353, -32'd2376, -32'd9030, 32'd2783},
{-32'd5934, 32'd4461, -32'd6659, -32'd553},
{-32'd11150, -32'd1005, -32'd10256, 32'd4773},
{-32'd7636, 32'd6511, -32'd10476, -32'd1375},
{-32'd4448, 32'd5857, -32'd1416, 32'd4305},
{32'd1304, -32'd11105, 32'd9620, -32'd18136},
{32'd3997, -32'd3149, -32'd9087, 32'd5200},
{-32'd424, 32'd7742, -32'd8780, -32'd9514},
{32'd1368, 32'd3324, -32'd7144, 32'd8165},
{-32'd938, -32'd4473, -32'd16611, -32'd775}
},
{{-32'd161, -32'd11180, -32'd6725, -32'd1592},
{-32'd2265, -32'd2594, -32'd7379, -32'd7434},
{-32'd6635, -32'd14675, -32'd2269, -32'd4369},
{32'd4757, 32'd7551, -32'd2901, 32'd7457},
{32'd21379, 32'd570, -32'd5714, -32'd3039},
{32'd9139, 32'd14438, -32'd2288, -32'd5539},
{32'd2062, -32'd7244, 32'd9321, 32'd4428},
{-32'd10519, 32'd1590, 32'd9169, 32'd5420},
{-32'd5237, 32'd4220, 32'd8444, 32'd10145},
{32'd7825, 32'd165, 32'd14586, 32'd7098},
{32'd6412, -32'd330, -32'd6507, -32'd843},
{32'd3298, 32'd10722, 32'd2304, -32'd9145},
{32'd1146, 32'd7156, 32'd3949, 32'd1199},
{-32'd13953, -32'd3116, -32'd7887, -32'd3064},
{-32'd14880, 32'd727, -32'd8296, 32'd6465},
{-32'd1802, 32'd9139, -32'd6206, -32'd6213},
{32'd10105, -32'd1144, 32'd2571, 32'd7786},
{-32'd397, -32'd2232, -32'd8463, 32'd3487},
{32'd12476, -32'd10635, -32'd6213, -32'd7332},
{-32'd3097, -32'd6946, -32'd13025, 32'd3989},
{-32'd6958, 32'd4046, -32'd10168, 32'd3069},
{-32'd12662, -32'd5664, -32'd12662, -32'd14393},
{32'd323, 32'd4011, -32'd7516, 32'd1541},
{32'd2697, -32'd4592, -32'd9905, 32'd1067},
{32'd5727, 32'd1107, 32'd5813, -32'd7915},
{-32'd3521, -32'd5328, -32'd11426, -32'd3197},
{-32'd9178, 32'd4096, -32'd6628, 32'd8546},
{32'd6836, 32'd8576, 32'd9899, 32'd3002},
{32'd2116, -32'd101, -32'd10400, 32'd5503},
{-32'd17247, -32'd18737, 32'd13810, 32'd7433},
{32'd3650, -32'd9395, -32'd15946, 32'd2214},
{-32'd4550, -32'd349, -32'd8650, -32'd8957},
{32'd18349, -32'd5245, 32'd11187, -32'd3985},
{-32'd7498, 32'd2447, -32'd4096, -32'd8495},
{32'd9044, 32'd4999, 32'd11892, 32'd7225},
{-32'd611, -32'd1482, -32'd104, 32'd5630},
{-32'd1117, -32'd521, -32'd2396, 32'd1385},
{-32'd7318, 32'd9009, 32'd4694, -32'd10697},
{-32'd5528, 32'd5639, 32'd4577, -32'd10610},
{-32'd18410, -32'd2283, 32'd5611, -32'd8928},
{-32'd651, 32'd11171, -32'd802, -32'd7168},
{32'd9011, -32'd4947, 32'd8685, 32'd15425},
{-32'd7122, 32'd280, 32'd5429, -32'd14075},
{-32'd12439, 32'd4963, -32'd8763, -32'd4052},
{32'd1056, -32'd3217, 32'd3185, 32'd249},
{-32'd14652, 32'd20902, 32'd1854, -32'd12718},
{-32'd4940, 32'd12091, -32'd2860, -32'd3681},
{32'd3532, 32'd7665, 32'd371, 32'd2987},
{-32'd2404, -32'd990, 32'd10954, -32'd6028},
{32'd2357, 32'd2212, 32'd4959, 32'd859},
{-32'd10518, -32'd15714, 32'd3428, 32'd1757},
{-32'd7242, 32'd7233, 32'd5887, -32'd16380},
{-32'd2911, 32'd10896, -32'd2251, -32'd3812},
{32'd11370, -32'd21858, -32'd6167, 32'd7873},
{32'd11598, 32'd3650, 32'd8241, 32'd786},
{-32'd6648, -32'd11156, -32'd13208, 32'd590},
{-32'd1283, 32'd659, -32'd1334, 32'd683},
{-32'd9274, -32'd15234, -32'd14936, -32'd2091},
{-32'd7474, 32'd1994, -32'd17670, -32'd8231},
{32'd1516, -32'd9160, -32'd7606, 32'd3882},
{32'd10535, 32'd8378, -32'd18779, 32'd9359},
{32'd3175, -32'd2565, 32'd8628, -32'd13446},
{-32'd9384, -32'd6227, -32'd16694, 32'd6665},
{-32'd4972, -32'd6855, -32'd2649, -32'd2262},
{32'd16727, -32'd1709, -32'd12772, -32'd13331},
{32'd1942, 32'd3763, 32'd8617, 32'd582},
{-32'd1364, 32'd3646, -32'd15077, -32'd5609},
{-32'd8223, 32'd15245, -32'd1987, -32'd799},
{32'd3565, -32'd2888, 32'd1995, -32'd2678},
{32'd4363, 32'd5523, -32'd1888, 32'd4354},
{-32'd599, -32'd4827, 32'd3938, 32'd12811},
{32'd13640, -32'd242, -32'd2298, 32'd2090},
{32'd8809, -32'd19418, -32'd5290, -32'd6690},
{32'd403, -32'd13588, -32'd3475, -32'd168},
{32'd10718, 32'd1200, -32'd263, 32'd6978},
{-32'd9826, -32'd5500, 32'd8058, -32'd2179},
{-32'd11516, -32'd3757, 32'd4661, -32'd8805},
{32'd4230, 32'd13723, -32'd2973, 32'd14909},
{32'd8283, 32'd3265, 32'd9055, 32'd5313},
{32'd1865, -32'd11320, 32'd6423, 32'd3085},
{32'd13199, 32'd2271, -32'd4981, -32'd10716},
{32'd1989, -32'd11435, 32'd10549, -32'd6454},
{-32'd1525, -32'd8595, -32'd7531, -32'd6544},
{32'd3304, -32'd2354, -32'd2503, -32'd6767},
{32'd9057, -32'd15489, 32'd1294, -32'd10412},
{32'd5960, -32'd5440, -32'd2130, -32'd2050},
{32'd487, -32'd5059, 32'd4181, -32'd10068},
{32'd3605, -32'd12942, -32'd15728, 32'd3149},
{-32'd18983, -32'd6835, -32'd369, 32'd7458},
{32'd6698, -32'd4778, -32'd5512, -32'd1960},
{32'd4485, 32'd221, 32'd11280, -32'd2443},
{32'd1495, -32'd2574, -32'd5257, -32'd9865},
{-32'd9275, -32'd7572, 32'd12383, -32'd1826},
{32'd7720, 32'd3734, 32'd2993, -32'd6579},
{-32'd9292, -32'd448, -32'd5959, 32'd2929},
{32'd11883, -32'd7856, -32'd6459, -32'd9299},
{32'd2204, -32'd5363, 32'd12486, -32'd1214},
{-32'd9036, 32'd4433, 32'd6617, 32'd12154},
{32'd9725, 32'd8005, 32'd7021, 32'd5465},
{32'd20088, -32'd1080, 32'd25733, 32'd7376},
{-32'd2484, 32'd10206, -32'd234, -32'd8749},
{-32'd6948, -32'd6606, 32'd4735, 32'd1509},
{-32'd1563, -32'd11377, 32'd988, -32'd10211},
{32'd16358, 32'd11722, -32'd12094, 32'd3403},
{-32'd7518, 32'd4327, -32'd8441, -32'd3463},
{32'd329, -32'd1937, 32'd2658, 32'd1759},
{-32'd8840, 32'd4993, -32'd81, 32'd2791},
{-32'd9869, 32'd6652, -32'd6637, -32'd15003},
{32'd11399, 32'd5964, 32'd15646, 32'd2354},
{-32'd3866, 32'd4350, -32'd15089, 32'd7734},
{-32'd493, -32'd17885, 32'd8422, -32'd7271},
{-32'd1642, -32'd12897, 32'd7890, 32'd2297},
{-32'd2913, 32'd928, 32'd3946, 32'd52},
{32'd11832, 32'd8143, 32'd7081, -32'd6461},
{-32'd3299, -32'd5161, 32'd1411, -32'd8066},
{-32'd7295, 32'd13704, -32'd362, 32'd5314},
{32'd7491, -32'd3547, 32'd1640, -32'd4262},
{-32'd8565, 32'd4585, 32'd5754, -32'd13233},
{32'd4143, -32'd10175, -32'd7974, 32'd6453},
{32'd2109, 32'd2839, 32'd2874, -32'd2556},
{32'd3687, -32'd529, 32'd1290, -32'd13036},
{-32'd2823, -32'd4036, -32'd8092, -32'd1665},
{32'd909, 32'd16793, 32'd2244, -32'd8266},
{-32'd2235, -32'd55, -32'd7076, 32'd11590},
{32'd14852, -32'd18217, -32'd5169, 32'd7304},
{-32'd6697, 32'd6401, 32'd5847, 32'd12239},
{-32'd242, -32'd7353, -32'd2425, 32'd4839},
{-32'd23565, -32'd1024, 32'd1548, 32'd1444},
{-32'd18812, -32'd3781, 32'd1094, 32'd2044},
{-32'd1669, -32'd890, -32'd5246, 32'd15568},
{32'd10684, -32'd4482, 32'd1245, 32'd4451},
{-32'd5964, 32'd2143, 32'd2952, -32'd3539},
{-32'd8927, -32'd504, -32'd15646, -32'd7117},
{32'd9536, -32'd2462, 32'd7820, -32'd6295},
{-32'd700, -32'd2176, 32'd10922, 32'd9671},
{-32'd160, -32'd23485, -32'd4517, 32'd4837},
{32'd506, 32'd1221, 32'd9086, 32'd6414},
{32'd4618, 32'd12318, -32'd3981, 32'd1826},
{32'd6880, 32'd862, -32'd5464, 32'd5725},
{-32'd8668, 32'd8838, -32'd1280, -32'd1490},
{-32'd2229, -32'd5812, 32'd5472, 32'd2431},
{32'd4153, -32'd4457, 32'd6801, 32'd4671},
{-32'd639, 32'd7574, -32'd13346, -32'd5461},
{32'd14040, -32'd6985, -32'd7822, 32'd855},
{32'd2204, -32'd1281, 32'd3210, 32'd723},
{-32'd6275, 32'd7087, 32'd16755, -32'd9594},
{-32'd10022, -32'd5737, -32'd6065, -32'd4712},
{32'd8644, -32'd16788, -32'd7200, -32'd3569},
{-32'd1851, 32'd5331, 32'd7690, -32'd905},
{-32'd7754, -32'd4980, -32'd12052, -32'd3042},
{32'd5920, 32'd2592, -32'd2813, -32'd1394},
{32'd1966, 32'd5242, 32'd2422, -32'd4592},
{-32'd2329, 32'd8363, -32'd4872, -32'd12288},
{32'd1272, 32'd4046, 32'd4298, 32'd1860},
{32'd5334, 32'd2032, -32'd7071, 32'd2730},
{-32'd10074, 32'd2274, 32'd5080, 32'd13512},
{32'd127, 32'd11615, -32'd8339, 32'd515},
{32'd13223, 32'd5370, 32'd300, -32'd3714},
{-32'd1682, 32'd8717, -32'd10971, -32'd3084},
{32'd6590, -32'd9304, 32'd14938, 32'd1795},
{32'd6490, 32'd4625, 32'd2381, 32'd910},
{-32'd665, -32'd2495, 32'd13179, 32'd3007},
{32'd7064, -32'd250, -32'd5768, -32'd812},
{32'd2040, -32'd5946, 32'd8049, -32'd3888},
{-32'd7994, 32'd12285, 32'd5024, -32'd1925},
{-32'd6144, -32'd3111, -32'd10790, -32'd1060},
{32'd7614, 32'd4196, -32'd4725, 32'd1807},
{-32'd19017, 32'd1443, -32'd3961, 32'd4415},
{32'd10751, 32'd3495, 32'd5441, -32'd20033},
{32'd1612, 32'd308, -32'd14163, -32'd2343},
{32'd2099, -32'd1615, 32'd6805, 32'd2557},
{-32'd10766, -32'd412, 32'd7669, 32'd9163},
{32'd2178, 32'd9751, 32'd12189, 32'd9327},
{-32'd5186, 32'd2834, 32'd615, 32'd2232},
{-32'd13917, 32'd367, -32'd12312, 32'd8171},
{32'd1575, -32'd5264, -32'd1707, -32'd10479},
{-32'd2348, 32'd5098, -32'd8748, -32'd1693},
{-32'd13177, -32'd807, 32'd4821, 32'd8282},
{-32'd15259, -32'd6372, -32'd2267, 32'd4221},
{-32'd2654, -32'd2764, -32'd8028, -32'd5956},
{-32'd6815, 32'd1837, -32'd903, 32'd534},
{-32'd2433, 32'd3739, -32'd1330, -32'd494},
{-32'd2505, 32'd14334, -32'd16289, -32'd10209},
{32'd4035, 32'd70, -32'd10222, 32'd3031},
{32'd1585, 32'd1895, -32'd9945, -32'd4636},
{32'd11096, -32'd579, -32'd697, 32'd5105},
{32'd4197, 32'd1731, 32'd7883, 32'd12722},
{-32'd6741, -32'd6072, 32'd14955, 32'd5668},
{-32'd9100, -32'd3427, -32'd2939, 32'd3824},
{32'd3385, -32'd4958, -32'd4725, 32'd7684},
{-32'd1725, 32'd1208, -32'd5592, 32'd3417},
{-32'd928, -32'd3641, -32'd968, 32'd1848},
{-32'd18974, -32'd1632, -32'd16742, -32'd7351},
{-32'd15695, 32'd7370, 32'd8560, 32'd423},
{32'd2529, -32'd7519, 32'd8216, 32'd12851},
{-32'd5603, -32'd3717, -32'd239, 32'd743},
{32'd7909, 32'd14960, -32'd8931, 32'd2856},
{32'd1289, -32'd4507, -32'd1959, 32'd1189},
{-32'd1312, -32'd6697, 32'd4258, 32'd5711},
{32'd18195, 32'd7294, 32'd5869, -32'd5813},
{-32'd4102, -32'd5098, -32'd12049, -32'd4619},
{32'd8069, 32'd2171, 32'd6934, -32'd10039},
{32'd15460, 32'd284, -32'd3559, -32'd3665},
{32'd645, 32'd5739, 32'd19272, 32'd3829},
{-32'd9151, -32'd12685, -32'd6517, -32'd15316},
{32'd13163, 32'd11980, 32'd2603, 32'd4328},
{-32'd14242, 32'd1063, -32'd583, 32'd1159},
{-32'd10857, 32'd6729, -32'd1899, -32'd5569},
{32'd9645, 32'd5449, -32'd2905, 32'd8579},
{-32'd2896, 32'd9809, 32'd6438, -32'd5178},
{32'd14423, 32'd128, 32'd5606, -32'd14463},
{-32'd3055, 32'd5922, 32'd4088, -32'd3363},
{-32'd659, -32'd14527, -32'd2057, 32'd5407},
{-32'd8222, 32'd6193, 32'd6748, -32'd6926},
{-32'd9725, -32'd11307, -32'd3933, -32'd16352},
{32'd12400, 32'd2338, -32'd13161, 32'd4523},
{32'd3472, -32'd6610, -32'd3938, 32'd7205},
{-32'd6429, 32'd5552, -32'd5785, 32'd2167},
{-32'd231, 32'd3128, 32'd1908, 32'd6819},
{32'd848, 32'd3165, -32'd2458, 32'd11522},
{-32'd15529, 32'd2014, 32'd122, 32'd2709},
{32'd10479, 32'd6132, -32'd7142, 32'd8812},
{-32'd1898, -32'd5319, -32'd1027, 32'd10744},
{32'd9552, 32'd3774, -32'd7900, -32'd3608},
{32'd1848, 32'd9283, -32'd14001, -32'd1355},
{32'd4579, 32'd14065, 32'd8408, -32'd15574},
{-32'd4999, 32'd3651, 32'd5216, -32'd2327},
{32'd1590, -32'd10535, -32'd4866, -32'd1393},
{-32'd9288, -32'd7842, 32'd1355, 32'd6785},
{-32'd7732, 32'd14777, 32'd7259, -32'd2453},
{-32'd12656, 32'd1786, 32'd1567, 32'd9377},
{-32'd4248, -32'd6391, 32'd2708, -32'd4983},
{32'd10493, -32'd53, -32'd913, 32'd9546},
{32'd14136, -32'd8930, 32'd14333, 32'd3412},
{32'd250, 32'd5442, -32'd6502, -32'd11527},
{-32'd10741, -32'd19634, -32'd368, 32'd524},
{32'd659, 32'd10561, -32'd5306, 32'd3643},
{-32'd11920, 32'd18411, 32'd1825, -32'd857},
{-32'd1238, 32'd10436, 32'd3320, 32'd2247},
{32'd1235, -32'd1533, 32'd2712, 32'd3618},
{-32'd5757, -32'd10828, 32'd3360, -32'd1824},
{-32'd3141, 32'd7618, -32'd5661, -32'd4589},
{32'd308, -32'd6366, -32'd13997, -32'd2527},
{-32'd13984, -32'd20364, 32'd4722, -32'd2405},
{32'd6981, 32'd3285, 32'd12863, 32'd3500},
{32'd2149, -32'd8083, 32'd6248, 32'd10053},
{32'd972, 32'd735, 32'd8317, -32'd3648},
{32'd9654, -32'd5879, -32'd4296, -32'd5048},
{32'd6014, -32'd447, -32'd1716, -32'd109},
{-32'd443, 32'd74, -32'd4981, -32'd6162},
{32'd8496, -32'd160, -32'd3861, 32'd3968},
{32'd7920, 32'd11157, 32'd16434, -32'd2247},
{32'd27779, 32'd9915, 32'd13966, 32'd3529},
{-32'd1412, 32'd20622, -32'd8908, -32'd1921},
{-32'd7493, -32'd1033, -32'd4734, -32'd11499},
{-32'd14242, 32'd5889, 32'd10525, 32'd3333},
{32'd3746, -32'd2144, -32'd6006, -32'd2723},
{32'd9910, -32'd14476, 32'd8240, -32'd3544},
{32'd5301, -32'd9975, -32'd1214, -32'd5865},
{32'd1684, -32'd2338, 32'd17585, -32'd5638},
{-32'd2543, 32'd2522, -32'd3729, 32'd6308},
{32'd4803, 32'd788, 32'd1675, 32'd6467},
{32'd1822, 32'd12554, -32'd5086, 32'd1228},
{-32'd9907, -32'd3175, 32'd3991, 32'd515},
{-32'd512, 32'd509, 32'd332, -32'd19839},
{32'd8702, -32'd9066, -32'd594, -32'd2153},
{32'd7023, -32'd2759, 32'd77, 32'd14333},
{32'd12220, -32'd4957, -32'd5046, -32'd2835},
{-32'd4190, -32'd7886, -32'd12467, 32'd1152},
{32'd2064, 32'd13901, -32'd7587, -32'd1518},
{32'd12568, 32'd2908, 32'd8491, 32'd1952},
{32'd5843, 32'd8547, 32'd8806, 32'd787},
{-32'd3154, -32'd537, -32'd14241, 32'd4404},
{-32'd2826, 32'd4924, 32'd11604, 32'd708},
{32'd11461, -32'd24, 32'd7597, -32'd13391},
{-32'd4370, -32'd6415, -32'd6978, 32'd4616},
{32'd10531, 32'd5082, 32'd13601, 32'd7889},
{-32'd9054, 32'd10480, 32'd9105, -32'd5262},
{32'd1370, -32'd1502, -32'd15460, -32'd3041},
{-32'd4050, 32'd5915, -32'd4981, -32'd3369},
{32'd7640, -32'd15531, 32'd3225, 32'd4987},
{-32'd19241, -32'd4416, 32'd7562, 32'd1952},
{32'd7643, -32'd5829, 32'd2299, 32'd14653},
{-32'd931, 32'd6876, -32'd175, 32'd2679},
{-32'd3394, 32'd5494, -32'd2998, -32'd2214},
{-32'd110, 32'd2600, -32'd13662, -32'd5922},
{32'd4432, -32'd15094, 32'd8285, 32'd5135},
{32'd11995, -32'd8205, 32'd9279, -32'd13131},
{32'd6106, 32'd5210, 32'd897, -32'd7112},
{-32'd20391, -32'd9802, -32'd1359, -32'd426},
{32'd4927, -32'd6846, 32'd7304, 32'd5687},
{32'd2022, -32'd6726, 32'd10786, 32'd5209},
{-32'd11451, -32'd20635, -32'd5087, -32'd2463},
{-32'd3354, 32'd6441, 32'd8143, -32'd4890},
{-32'd2687, -32'd13409, -32'd3663, 32'd9654},
{32'd1247, -32'd2376, 32'd2837, -32'd3016},
{-32'd510, -32'd5539, 32'd583, -32'd5808},
{32'd7667, 32'd1770, 32'd7749, -32'd6881},
{-32'd1419, 32'd6138, 32'd10153, 32'd13023},
{32'd2505, -32'd6502, -32'd17845, -32'd3199}
}
};
